module SOMAMAISMAIS (A, B, S);
input [7:0] A;
input [3:0] B;
output reg [7:0] S;
always @(*)
begin
    if(A == 8'b00000000) begin
        if(B == 4'b0000) begin
            S = 8'b00000000;
        end
    end
    if(A == 8'b00000001) begin
        if(B == 4'b0000) begin
            S = 8'b00000001;
        end
    end
    if(A == 8'b00000010) begin
        if(B == 4'b0000) begin
            S = 8'b00000010;
        end
    end
    if(A == 8'b00000011) begin
        if(B == 4'b0000) begin
            S = 8'b00000011;
        end
    end
    if(A == 8'b00000100) begin
        if(B == 4'b0000) begin
            S = 8'b00000100;
        end
    end
    if(A == 8'b00000101) begin
        if(B == 4'b0000) begin
            S = 8'b00000101;
        end
    end
    if(A == 8'b00000110) begin
        if(B == 4'b0000) begin
            S = 8'b00000110;
        end
    end
    if(A == 8'b00000111) begin
        if(B == 4'b0000) begin
            S = 8'b00000111;
        end
    end
    if(A == 8'b00001000) begin
        if(B == 4'b0000) begin
            S = 8'b00001000;
        end
    end
    if(A == 8'b00001001) begin
        if(B == 4'b0000) begin
            S = 8'b00001001;
        end
    end
    if(A == 8'b00001010) begin
        if(B == 4'b0000) begin
            S = 8'b00001010;
        end
    end
    if(A == 8'b00001011) begin
        if(B == 4'b0000) begin
            S = 8'b00001011;
        end
    end
    if(A == 8'b00001100) begin
        if(B == 4'b0000) begin
            S = 8'b00001100;
        end
    end
    if(A == 8'b00001101) begin
        if(B == 4'b0000) begin
            S = 8'b00001101;
        end
    end
    if(A == 8'b00001110) begin
        if(B == 4'b0000) begin
            S = 8'b00001110;
        end
    end
    if(A == 8'b00001111) begin
        if(B == 4'b0000) begin
            S = 8'b00001111;
        end
    end
    if(A == 8'b00010000) begin
        if(B == 4'b0000) begin
            S = 8'b00010000;
        end
    end
    if(A == 8'b000010001) begin
        if(B == 4'b0000) begin
            S = 8'b000010001;
        end
    end
    if(A == 8'b000010010) begin
        if(B == 4'b0000) begin
            S = 8'b000010010;
        end
    end
    if(A == 8'b000010011) begin
        if(B == 4'b0000) begin
            S = 8'b000010011;
        end
    end
    if(A == 8'b000010100) begin
        if(B == 4'b0000) begin
            S = 8'b000010100;
        end
    end
    if(A == 8'b000010101) begin
        if(B == 4'b0000) begin
            S = 8'b000010101;
        end
    end
    if(A == 8'b000010110) begin
        if(B == 4'b0000) begin
            S = 8'b000010110;
        end
    end
    if(A == 8'b000010111) begin
        if(B == 4'b0000) begin
            S = 8'b000010111;
        end
    end
    if(A == 8'b00011000) begin
        if(B == 4'b0000) begin
            S = 8'b00011000;
        end
    end
    if(A == 8'b00011001) begin
        if(B == 4'b0000) begin
            S = 8'b00011001;
        end
    end
    if(A == 8'b00011010) begin
        if(B == 4'b0000) begin
            S = 8'b00011010;
        end
    end
    if(A == 8'b00011011) begin
        if(B == 4'b0000) begin
            S = 8'b00011011;
        end
    end
    if(A == 8'b00011100) begin
        if(B == 4'b0000) begin
            S = 8'b00011100;
        end
    end
    if(A == 8'b00011101) begin
        if(B == 4'b0000) begin
            S = 8'b00011101;
        end
    end
    if(A == 8'b00011110) begin
        if(B == 4'b0000) begin
            S = 8'b00011110;
        end
    end
    if(A == 8'b00011111) begin
        if(B == 4'b0000) begin
            S = 8'b00011111;
        end
    end
    if(A == 8'b00100000) begin
        if(B == 4'b0000) begin
            S = 8'b00100000;
        end
    end
    if(A == 8'b00100001) begin
        if(B == 4'b0000) begin
            S = 8'b00100001;
        end
    end
    if(A == 8'b00100010) begin
        if(B == 4'b0000) begin
            S = 8'b00100010;
        end
    end
    if(A == 8'b00100011) begin
        if(B == 4'b0000) begin
            S = 8'b00100011;
        end
    end
    if(A == 8'b00100100) begin
        if(B == 4'b0000) begin
            S = 8'b00100100;
        end
    end
    if(A == 8'b00100101) begin
        if(B == 4'b0000) begin
            S = 8'b00100101;
        end
    end
    if(A == 8'b00100110) begin
        if(B == 4'b0000) begin
            S = 8'b00100110;
        end
    end
    if(A == 8'b00100111) begin
        if(B == 4'b0000) begin
            S = 8'b00100111;
        end
    end
    if(A == 8'b00101000) begin
        if(B == 4'b0000) begin
            S = 8'b00101000;
        end
    end
    if(A == 8'b00101001) begin
        if(B == 4'b0000) begin
            S = 8'b00101001;
        end
    end
    if(A == 8'b00101010) begin
        if(B == 4'b0000) begin
            S = 8'b00101010;
        end
    end
    if(A == 8'b00101011) begin
        if(B == 4'b0000) begin
            S = 8'b00101011;
        end
    end
    if(A == 8'b00101100) begin
        if(B == 4'b0000) begin
            S = 8'b00101100;
        end
    end
    if(A == 8'b00101101) begin
        if(B == 4'b0000) begin
            S = 8'b00101101;
        end
    end
    if(A == 8'b00101110) begin
        if(B == 4'b0000) begin
            S = 8'b00101110;
        end
    end
    if(A == 8'b00101111) begin
        if(B == 4'b0000) begin
            S = 8'b00101111;
        end
    end
    if(A == 8'b00110000) begin
        if(B == 4'b0000) begin
            S = 8'b00110000;
        end
    end
    if(A == 8'b00110001) begin
        if(B == 4'b0000) begin
            S = 8'b00110001;
        end
    end
    if(A == 8'b00110010) begin
        if(B == 4'b0000) begin
            S = 8'b00110010;
        end
    end
    if(A == 8'b00110011) begin
        if(B == 4'b0000) begin
            S = 8'b00110011;
        end
    end
    if(A == 8'b00110100) begin
        if(B == 4'b0000) begin
            S = 8'b00110100;
        end
    end
    if(A == 8'b00110101) begin
        if(B == 4'b0000) begin
            S = 8'b00110101;
        end
    end
    if(A == 8'b00110110) begin
        if(B == 4'b0000) begin
            S = 8'b00110110;
        end
    end
    if(A == 8'b00110111) begin
        if(B == 4'b0000) begin
            S = 8'b00110111;
        end
    end
    if(A == 8'b00111000) begin
        if(B == 4'b0000) begin
            S = 8'b00111000;
        end
    end
    if(A == 8'b00111001) begin
        if(B == 4'b0000) begin
            S = 8'b00111001;
        end
    end
    if(A == 8'b00111010) begin
        if(B == 4'b0000) begin
            S = 8'b00111010;
        end
    end
    if(A == 8'b00111011) begin
        if(B == 4'b0000) begin
            S = 8'b00111011;
        end
    end
    if(A == 8'b00111100) begin
        if(B == 4'b0000) begin
            S = 8'b00111100;
        end
    end
    if(A == 8'b00111101) begin
        if(B == 4'b0000) begin
            S = 8'b00111101;
        end
    end
    if(A == 8'b00111110) begin
        if(B == 4'b0000) begin
            S = 8'b00111110;
        end
    end
    if(A == 8'b00111111) begin
        if(B == 4'b0000) begin
            S = 8'b00111111;
        end
    end
    if(A == 8'b01000000) begin
        if(B == 4'b0000) begin
            S = 8'b01000000;
        end
    end
    if(A == 8'b01000001) begin
        if(B == 4'b0000) begin
            S = 8'b01000001;
        end
    end
    if(A == 8'b01000010) begin
        if(B == 4'b0000) begin
            S = 8'b01000010;
        end
    end
    if(A == 8'b01000011) begin
        if(B == 4'b0000) begin
            S = 8'b01000011;
        end
    end
    if(A == 8'b01000100) begin
        if(B == 4'b0000) begin
            S = 8'b01000100;
        end
    end
    if(A == 8'b01000101) begin
        if(B == 4'b0000) begin
            S = 8'b01000101;
        end
    end
    if(A == 8'b01000110) begin
        if(B == 4'b0000) begin
            S = 8'b01000110;
        end
    end
    if(A == 8'b01000111) begin
        if(B == 4'b0000) begin
            S = 8'b01000111;
        end
    end
    if(A == 8'b01001000) begin
        if(B == 4'b0000) begin
            S = 8'b01001000;
        end
    end
    if(A == 8'b01001001) begin
        if(B == 4'b0000) begin
            S = 8'b01001001;
        end
    end
    if(A == 8'b01001010) begin
        if(B == 4'b0000) begin
            S = 8'b01001010;
        end
    end
    if(A == 8'b01001011) begin
        if(B == 4'b0000) begin
            S = 8'b01001011;
        end
    end
    if(A == 8'b01001100) begin
        if(B == 4'b0000) begin
            S = 8'b01001100;
        end
    end
    if(A == 8'b01001101) begin
        if(B == 4'b0000) begin
            S = 8'b01001101;
        end
    end
    if(A == 8'b01001110) begin
        if(B == 4'b0000) begin
            S = 8'b01001110;
        end
    end
    if(A == 8'b01001111) begin
        if(B == 4'b0000) begin
            S = 8'b01001111;
        end
    end
    if(A == 8'b01010000) begin
        if(B == 4'b0000) begin
            S = 8'b01010000;
        end
    end
    if(A == 8'b01010001) begin
        if(B == 4'b0000) begin
            S = 8'b01010001;
        end
    end
    if(A == 8'b01010010) begin
        if(B == 4'b0000) begin
            S = 8'b01010010;
        end
    end
    if(A == 8'b01010011) begin
        if(B == 4'b0000) begin
            S = 8'b01010011;
        end
    end
    if(A == 8'b01010100) begin
        if(B == 4'b0000) begin
            S = 8'b01010100;
        end
    end
    if(A == 8'b01010101) begin
        if(B == 4'b0000) begin
            S = 8'b01010101;
        end
    end
    if(A == 8'b01010110) begin
        if(B == 4'b0000) begin
            S = 8'b01010110;
        end
    end
    if(A == 8'b01010111) begin
        if(B == 4'b0000) begin
            S = 8'b01010111;
        end
    end
    if(A == 8'b01011000) begin
        if(B == 4'b0000) begin
            S = 8'b01011000;
        end
    end
    if(A == 8'b01011001) begin
        if(B == 4'b0000) begin
            S = 8'b01011001;
        end
    end
    if(A == 8'b01011010) begin
        if(B == 4'b0000) begin
            S = 8'b01011010;
        end
    end
    if(A == 8'b01011011) begin
        if(B == 4'b0000) begin
            S = 8'b01011011;
        end
    end
    if(A == 8'b01011100) begin
        if(B == 4'b0000) begin
            S = 8'b01011100;
        end
    end
    if(A == 8'b01011101) begin
        if(B == 4'b0000) begin
            S = 8'b01011101;
        end
    end
    if(A == 8'b01011110) begin
        if(B == 4'b0000) begin
            S = 8'b01011110;
        end
    end
    if(A == 8'b01011111) begin
        if(B == 4'b0000) begin
            S = 8'b01011111;
        end
    end
    if(A == 8'b01100000) begin
        if(B == 4'b0000) begin
            S = 8'b01100000;
        end
    end
    if(A == 8'b01100001) begin
        if(B == 4'b0000) begin
            S = 8'b01100001;
        end
    end
    if(A == 8'b01100010) begin
        if(B == 4'b0000) begin
            S = 8'b01100010;
        end
    end
    if(A == 8'b01100011) begin
        if(B == 4'b0000) begin
            S = 8'b01100011;
        end
    end
    if(A == 8'b00000000) begin
        if(B == 4'b0001) begin
            S = 8'b00000001;
        end
    end
    if(A == 8'b00000001) begin
        if(B == 4'b0001) begin
            S = 8'b00000010;
        end
    end
    if(A == 8'b00000010) begin
        if(B == 4'b0001) begin
            S = 8'b00000011;
        end
    end
    if(A == 8'b00000011) begin
        if(B == 4'b0001) begin
            S = 8'b00000100;
        end
    end
    if(A == 8'b00000100) begin
        if(B == 4'b0001) begin
            S = 8'b00000101;
        end
    end
    if(A == 8'b00000101) begin
        if(B == 4'b0001) begin
            S = 8'b00000110;
        end
    end
    if(A == 8'b00000110) begin
        if(B == 4'b0001) begin
            S = 8'b00000111;
        end
    end
    if(A == 8'b00000111) begin
        if(B == 4'b0001) begin
            S = 8'b00001000;
        end
    end
    if(A == 8'b00001000) begin
        if(B == 4'b0001) begin
            S = 8'b00001001;
        end
    end
    if(A == 8'b00001001) begin
        if(B == 4'b0001) begin
            S = 8'b00001010;
        end
    end
    if(A == 8'b00001010) begin
        if(B == 4'b0001) begin
            S = 8'b00001011;
        end
    end
    if(A == 8'b00001011) begin
        if(B == 4'b0001) begin
            S = 8'b00001100;
        end
    end
    if(A == 8'b00001100) begin
        if(B == 4'b0001) begin
            S = 8'b00001101;
        end
    end
    if(A == 8'b00001101) begin
        if(B == 4'b0001) begin
            S = 8'b00001110;
        end
    end
    if(A == 8'b00001110) begin
        if(B == 4'b0001) begin
            S = 8'b00001111;
        end
    end
    if(A == 8'b00001111) begin
        if(B == 4'b0001) begin
            S = 8'b00010000;
        end
    end
    if(A == 8'b00010000) begin
        if(B == 4'b0001) begin
            S = 8'b000010001;
        end
    end
    if(A == 8'b000010001) begin
        if(B == 4'b0001) begin
            S = 8'b000010010;
        end
    end
    if(A == 8'b000010010) begin
        if(B == 4'b0001) begin
            S = 8'b000010011;
        end
    end
    if(A == 8'b000010011) begin
        if(B == 4'b0001) begin
            S = 8'b000010100;
        end
    end
    if(A == 8'b000010100) begin
        if(B == 4'b0001) begin
            S = 8'b000010101;
        end
    end
    if(A == 8'b000010101) begin
        if(B == 4'b0001) begin
            S = 8'b000010110;
        end
    end
    if(A == 8'b000010110) begin
        if(B == 4'b0001) begin
            S = 8'b000010111;
        end
    end
    if(A == 8'b000010111) begin
        if(B == 4'b0001) begin
            S = 8'b00011000;
        end
    end
    if(A == 8'b00011000) begin
        if(B == 4'b0001) begin
            S = 8'b00011001;
        end
    end
    if(A == 8'b00011001) begin
        if(B == 4'b0001) begin
            S = 8'b00011010;
        end
    end
    if(A == 8'b00011010) begin
        if(B == 4'b0001) begin
            S = 8'b00011011;
        end
    end
    if(A == 8'b00011011) begin
        if(B == 4'b0001) begin
            S = 8'b00011100;
        end
    end
    if(A == 8'b00011100) begin
        if(B == 4'b0001) begin
            S = 8'b00011101;
        end
    end
    if(A == 8'b00011101) begin
        if(B == 4'b0001) begin
            S = 8'b00011110;
        end
    end
    if(A == 8'b00011110) begin
        if(B == 4'b0001) begin
            S = 8'b00011111;
        end
    end
    if(A == 8'b00011111) begin
        if(B == 4'b0001) begin
            S = 8'b00100000;
        end
    end
    if(A == 8'b00100000) begin
        if(B == 4'b0001) begin
            S = 8'b00100001;
        end
    end
    if(A == 8'b00100001) begin
        if(B == 4'b0001) begin
            S = 8'b00100010;
        end
    end
    if(A == 8'b00100010) begin
        if(B == 4'b0001) begin
            S = 8'b00100011;
        end
    end
    if(A == 8'b00100011) begin
        if(B == 4'b0001) begin
            S = 8'b00100100;
        end
    end
    if(A == 8'b00100100) begin
        if(B == 4'b0001) begin
            S = 8'b00100101;
        end
    end
    if(A == 8'b00100101) begin
        if(B == 4'b0001) begin
            S = 8'b00100110;
        end
    end
    if(A == 8'b00100110) begin
        if(B == 4'b0001) begin
            S = 8'b00100111;
        end
    end
    if(A == 8'b00100111) begin
        if(B == 4'b0001) begin
            S = 8'b00101000;
        end
    end
    if(A == 8'b00101000) begin
        if(B == 4'b0001) begin
            S = 8'b00101001;
        end
    end
    if(A == 8'b00101001) begin
        if(B == 4'b0001) begin
            S = 8'b00101010;
        end
    end
    if(A == 8'b00101010) begin
        if(B == 4'b0001) begin
            S = 8'b00101011;
        end
    end
    if(A == 8'b00101011) begin
        if(B == 4'b0001) begin
            S = 8'b00101100;
        end
    end
    if(A == 8'b00101100) begin
        if(B == 4'b0001) begin
            S = 8'b00101101;
        end
    end
    if(A == 8'b00101101) begin
        if(B == 4'b0001) begin
            S = 8'b00101110;
        end
    end
    if(A == 8'b00101110) begin
        if(B == 4'b0001) begin
            S = 8'b00101111;
        end
    end
    if(A == 8'b00101111) begin
        if(B == 4'b0001) begin
            S = 8'b00110000;
        end
    end
    if(A == 8'b00110000) begin
        if(B == 4'b0001) begin
            S = 8'b00110001;
        end
    end
    if(A == 8'b00110001) begin
        if(B == 4'b0001) begin
            S = 8'b00110010;
        end
    end
    if(A == 8'b00110010) begin
        if(B == 4'b0001) begin
            S = 8'b00110011;
        end
    end
    if(A == 8'b00110011) begin
        if(B == 4'b0001) begin
            S = 8'b00110100;
        end
    end
    if(A == 8'b00110100) begin
        if(B == 4'b0001) begin
            S = 8'b00110101;
        end
    end
    if(A == 8'b00110101) begin
        if(B == 4'b0001) begin
            S = 8'b00110110;
        end
    end
    if(A == 8'b00110110) begin
        if(B == 4'b0001) begin
            S = 8'b00110111;
        end
    end
    if(A == 8'b00110111) begin
        if(B == 4'b0001) begin
            S = 8'b00111000;
        end
    end
    if(A == 8'b00111000) begin
        if(B == 4'b0001) begin
            S = 8'b00111001;
        end
    end
    if(A == 8'b00111001) begin
        if(B == 4'b0001) begin
            S = 8'b00111010;
        end
    end
    if(A == 8'b00111010) begin
        if(B == 4'b0001) begin
            S = 8'b00111011;
        end
    end
    if(A == 8'b00111011) begin
        if(B == 4'b0001) begin
            S = 8'b00111100;
        end
    end
    if(A == 8'b00111100) begin
        if(B == 4'b0001) begin
            S = 8'b00111101;
        end
    end
    if(A == 8'b00111101) begin
        if(B == 4'b0001) begin
            S = 8'b00111110;
        end
    end
    if(A == 8'b00111110) begin
        if(B == 4'b0001) begin
            S = 8'b00111111;
        end
    end
    if(A == 8'b00111111) begin
        if(B == 4'b0001) begin
            S = 8'b01000000;
        end
    end
    if(A == 8'b01000000) begin
        if(B == 4'b0001) begin
            S = 8'b01000001;
        end
    end
    if(A == 8'b01000001) begin
        if(B == 4'b0001) begin
            S = 8'b01000010;
        end
    end
    if(A == 8'b01000010) begin
        if(B == 4'b0001) begin
            S = 8'b01000011;
        end
    end
    if(A == 8'b01000011) begin
        if(B == 4'b0001) begin
            S = 8'b01000100;
        end
    end
    if(A == 8'b01000100) begin
        if(B == 4'b0001) begin
            S = 8'b01000101;
        end
    end
    if(A == 8'b01000101) begin
        if(B == 4'b0001) begin
            S = 8'b01000110;
        end
    end
    if(A == 8'b01000110) begin
        if(B == 4'b0001) begin
            S = 8'b01000111;
        end
    end
    if(A == 8'b01000111) begin
        if(B == 4'b0001) begin
            S = 8'b01001000;
        end
    end
    if(A == 8'b01001000) begin
        if(B == 4'b0001) begin
            S = 8'b01001001;
        end
    end
    if(A == 8'b01001001) begin
        if(B == 4'b0001) begin
            S = 8'b01001010;
        end
    end
    if(A == 8'b01001010) begin
        if(B == 4'b0001) begin
            S = 8'b01001011;
        end
    end
    if(A == 8'b01001011) begin
        if(B == 4'b0001) begin
            S = 8'b01001100;
        end
    end
    if(A == 8'b01001100) begin
        if(B == 4'b0001) begin
            S = 8'b01001101;
        end
    end
    if(A == 8'b01001101) begin
        if(B == 4'b0001) begin
            S = 8'b01001110;
        end
    end
    if(A == 8'b01001110) begin
        if(B == 4'b0001) begin
            S = 8'b01001111;
        end
    end
    if(A == 8'b01001111) begin
        if(B == 4'b0001) begin
            S = 8'b01010000;
        end
    end
    if(A == 8'b01010000) begin
        if(B == 4'b0001) begin
            S = 8'b01010001;
        end
    end
    if(A == 8'b01010001) begin
        if(B == 4'b0001) begin
            S = 8'b01010010;
        end
    end
    if(A == 8'b01010010) begin
        if(B == 4'b0001) begin
            S = 8'b01010011;
        end
    end
    if(A == 8'b01010011) begin
        if(B == 4'b0001) begin
            S = 8'b01010100;
        end
    end
    if(A == 8'b01010100) begin
        if(B == 4'b0001) begin
            S = 8'b01010101;
        end
    end
    if(A == 8'b01010101) begin
        if(B == 4'b0001) begin
            S = 8'b01010110;
        end
    end
    if(A == 8'b01010110) begin
        if(B == 4'b0001) begin
            S = 8'b01010111;
        end
    end
    if(A == 8'b01010111) begin
        if(B == 4'b0001) begin
            S = 8'b01011000;
        end
    end
    if(A == 8'b01011000) begin
        if(B == 4'b0001) begin
            S = 8'b01011001;
        end
    end
    if(A == 8'b01011001) begin
        if(B == 4'b0001) begin
            S = 8'b01011010;
        end
    end
    if(A == 8'b01011010) begin
        if(B == 4'b0001) begin
            S = 8'b01011011;
        end
    end
    if(A == 8'b01011011) begin
        if(B == 4'b0001) begin
            S = 8'b01011100;
        end
    end
    if(A == 8'b01011100) begin
        if(B == 4'b0001) begin
            S = 8'b01011101;
        end
    end
    if(A == 8'b01011101) begin
        if(B == 4'b0001) begin
            S = 8'b01011110;
        end
    end
    if(A == 8'b01011110) begin
        if(B == 4'b0001) begin
            S = 8'b01011111;
        end
    end
    if(A == 8'b01011111) begin
        if(B == 4'b0001) begin
            S = 8'b01100000;
        end
    end
    if(A == 8'b01100000) begin
        if(B == 4'b0001) begin
            S = 8'b01100001;
        end
    end
    if(A == 8'b01100001) begin
        if(B == 4'b0001) begin
            S = 8'b01100010;
        end
    end
    if(A == 8'b01100010) begin
        if(B == 4'b0001) begin
            S = 8'b01100011;
        end
    end
    if(A == 8'b00000000) begin
        if(B == 4'b0010) begin
            S = 8'b00000010;
        end
    end
    if(A == 8'b00000001) begin
        if(B == 4'b0010) begin
            S = 8'b00000011;
        end
    end
    if(A == 8'b00000010) begin
        if(B == 4'b0010) begin
            S = 8'b00000100;
        end
    end
    if(A == 8'b00000011) begin
        if(B == 4'b0010) begin
            S = 8'b00000101;
        end
    end
    if(A == 8'b00000100) begin
        if(B == 4'b0010) begin
            S = 8'b00000110;
        end
    end
    if(A == 8'b00000101) begin
        if(B == 4'b0010) begin
            S = 8'b00000111;
        end
    end
    if(A == 8'b00000110) begin
        if(B == 4'b0010) begin
            S = 8'b00001000;
        end
    end
    if(A == 8'b00000111) begin
        if(B == 4'b0010) begin
            S = 8'b00001001;
        end
    end
    if(A == 8'b00001000) begin
        if(B == 4'b0010) begin
            S = 8'b00001010;
        end
    end
    if(A == 8'b00001001) begin
        if(B == 4'b0010) begin
            S = 8'b00001011;
        end
    end
    if(A == 8'b00001010) begin
        if(B == 4'b0010) begin
            S = 8'b00001100;
        end
    end
    if(A == 8'b00001011) begin
        if(B == 4'b0010) begin
            S = 8'b00001101;
        end
    end
    if(A == 8'b00001100) begin
        if(B == 4'b0010) begin
            S = 8'b00001110;
        end
    end
    if(A == 8'b00001101) begin
        if(B == 4'b0010) begin
            S = 8'b00001111;
        end
    end
    if(A == 8'b00001110) begin
        if(B == 4'b0010) begin
            S = 8'b00010000;
        end
    end
    if(A == 8'b00001111) begin
        if(B == 4'b0010) begin
            S = 8'b000010001;
        end
    end
    if(A == 8'b00010000) begin
        if(B == 4'b0010) begin
            S = 8'b000010010;
        end
    end
    if(A == 8'b000010001) begin
        if(B == 4'b0010) begin
            S = 8'b000010011;
        end
    end
    if(A == 8'b000010010) begin
        if(B == 4'b0010) begin
            S = 8'b000010100;
        end
    end
    if(A == 8'b000010011) begin
        if(B == 4'b0010) begin
            S = 8'b000010101;
        end
    end
    if(A == 8'b000010100) begin
        if(B == 4'b0010) begin
            S = 8'b000010110;
        end
    end
    if(A == 8'b000010101) begin
        if(B == 4'b0010) begin
            S = 8'b000010111;
        end
    end
    if(A == 8'b000010110) begin
        if(B == 4'b0010) begin
            S = 8'b00011000;
        end
    end
    if(A == 8'b000010111) begin
        if(B == 4'b0010) begin
            S = 8'b00011001;
        end
    end
    if(A == 8'b00011000) begin
        if(B == 4'b0010) begin
            S = 8'b00011010;
        end
    end
    if(A == 8'b00011001) begin
        if(B == 4'b0010) begin
            S = 8'b00011011;
        end
    end
    if(A == 8'b00011010) begin
        if(B == 4'b0010) begin
            S = 8'b00011100;
        end
    end
    if(A == 8'b00011011) begin
        if(B == 4'b0010) begin
            S = 8'b00011101;
        end
    end
    if(A == 8'b00011100) begin
        if(B == 4'b0010) begin
            S = 8'b00011110;
        end
    end
    if(A == 8'b00011101) begin
        if(B == 4'b0010) begin
            S = 8'b00011111;
        end
    end
    if(A == 8'b00011110) begin
        if(B == 4'b0010) begin
            S = 8'b00100000;
        end
    end
    if(A == 8'b00011111) begin
        if(B == 4'b0010) begin
            S = 8'b00100001;
        end
    end
    if(A == 8'b00100000) begin
        if(B == 4'b0010) begin
            S = 8'b00100010;
        end
    end
    if(A == 8'b00100001) begin
        if(B == 4'b0010) begin
            S = 8'b00100011;
        end
    end
    if(A == 8'b00100010) begin
        if(B == 4'b0010) begin
            S = 8'b00100100;
        end
    end
    if(A == 8'b00100011) begin
        if(B == 4'b0010) begin
            S = 8'b00100101;
        end
    end
    if(A == 8'b00100100) begin
        if(B == 4'b0010) begin
            S = 8'b00100110;
        end
    end
    if(A == 8'b00100101) begin
        if(B == 4'b0010) begin
            S = 8'b00100111;
        end
    end
    if(A == 8'b00100110) begin
        if(B == 4'b0010) begin
            S = 8'b00101000;
        end
    end
    if(A == 8'b00100111) begin
        if(B == 4'b0010) begin
            S = 8'b00101001;
        end
    end
    if(A == 8'b00101000) begin
        if(B == 4'b0010) begin
            S = 8'b00101010;
        end
    end
    if(A == 8'b00101001) begin
        if(B == 4'b0010) begin
            S = 8'b00101011;
        end
    end
    if(A == 8'b00101010) begin
        if(B == 4'b0010) begin
            S = 8'b00101100;
        end
    end
    if(A == 8'b00101011) begin
        if(B == 4'b0010) begin
            S = 8'b00101101;
        end
    end
    if(A == 8'b00101100) begin
        if(B == 4'b0010) begin
            S = 8'b00101110;
        end
    end
    if(A == 8'b00101101) begin
        if(B == 4'b0010) begin
            S = 8'b00101111;
        end
    end
    if(A == 8'b00101110) begin
        if(B == 4'b0010) begin
            S = 8'b00110000;
        end
    end
    if(A == 8'b00101111) begin
        if(B == 4'b0010) begin
            S = 8'b00110001;
        end
    end
    if(A == 8'b00110000) begin
        if(B == 4'b0010) begin
            S = 8'b00110010;
        end
    end
    if(A == 8'b00110001) begin
        if(B == 4'b0010) begin
            S = 8'b00110011;
        end
    end
    if(A == 8'b00110010) begin
        if(B == 4'b0010) begin
            S = 8'b00110100;
        end
    end
    if(A == 8'b00110011) begin
        if(B == 4'b0010) begin
            S = 8'b00110101;
        end
    end
    if(A == 8'b00110100) begin
        if(B == 4'b0010) begin
            S = 8'b00110110;
        end
    end
    if(A == 8'b00110101) begin
        if(B == 4'b0010) begin
            S = 8'b00110111;
        end
    end
    if(A == 8'b00110110) begin
        if(B == 4'b0010) begin
            S = 8'b00111000;
        end
    end
    if(A == 8'b00110111) begin
        if(B == 4'b0010) begin
            S = 8'b00111001;
        end
    end
    if(A == 8'b00111000) begin
        if(B == 4'b0010) begin
            S = 8'b00111010;
        end
    end
    if(A == 8'b00111001) begin
        if(B == 4'b0010) begin
            S = 8'b00111011;
        end
    end
    if(A == 8'b00111010) begin
        if(B == 4'b0010) begin
            S = 8'b00111100;
        end
    end
    if(A == 8'b00111011) begin
        if(B == 4'b0010) begin
            S = 8'b00111101;
        end
    end
    if(A == 8'b00111100) begin
        if(B == 4'b0010) begin
            S = 8'b00111110;
        end
    end
    if(A == 8'b00111101) begin
        if(B == 4'b0010) begin
            S = 8'b00111111;
        end
    end
    if(A == 8'b00111110) begin
        if(B == 4'b0010) begin
            S = 8'b01000000;
        end
    end
    if(A == 8'b00111111) begin
        if(B == 4'b0010) begin
            S = 8'b01000001;
        end
    end
    if(A == 8'b01000000) begin
        if(B == 4'b0010) begin
            S = 8'b01000010;
        end
    end
    if(A == 8'b01000001) begin
        if(B == 4'b0010) begin
            S = 8'b01000011;
        end
    end
    if(A == 8'b01000010) begin
        if(B == 4'b0010) begin
            S = 8'b01000100;
        end
    end
    if(A == 8'b01000011) begin
        if(B == 4'b0010) begin
            S = 8'b01000101;
        end
    end
    if(A == 8'b01000100) begin
        if(B == 4'b0010) begin
            S = 8'b01000110;
        end
    end
    if(A == 8'b01000101) begin
        if(B == 4'b0010) begin
            S = 8'b01000111;
        end
    end
    if(A == 8'b01000110) begin
        if(B == 4'b0010) begin
            S = 8'b01001000;
        end
    end
    if(A == 8'b01000111) begin
        if(B == 4'b0010) begin
            S = 8'b01001001;
        end
    end
    if(A == 8'b01001000) begin
        if(B == 4'b0010) begin
            S = 8'b01001010;
        end
    end
    if(A == 8'b01001001) begin
        if(B == 4'b0010) begin
            S = 8'b01001011;
        end
    end
    if(A == 8'b01001010) begin
        if(B == 4'b0010) begin
            S = 8'b01001100;
        end
    end
    if(A == 8'b01001011) begin
        if(B == 4'b0010) begin
            S = 8'b01001101;
        end
    end
    if(A == 8'b01001100) begin
        if(B == 4'b0010) begin
            S = 8'b01001110;
        end
    end
    if(A == 8'b01001101) begin
        if(B == 4'b0010) begin
            S = 8'b01001111;
        end
    end
    if(A == 8'b01001110) begin
        if(B == 4'b0010) begin
            S = 8'b01010000;
        end
    end
    if(A == 8'b01001111) begin
        if(B == 4'b0010) begin
            S = 8'b01010001;
        end
    end
    if(A == 8'b01010000) begin
        if(B == 4'b0010) begin
            S = 8'b01010010;
        end
    end
    if(A == 8'b01010001) begin
        if(B == 4'b0010) begin
            S = 8'b01010011;
        end
    end
    if(A == 8'b01010010) begin
        if(B == 4'b0010) begin
            S = 8'b01010100;
        end
    end
    if(A == 8'b01010011) begin
        if(B == 4'b0010) begin
            S = 8'b01010101;
        end
    end
    if(A == 8'b01010100) begin
        if(B == 4'b0010) begin
            S = 8'b01010110;
        end
    end
    if(A == 8'b01010101) begin
        if(B == 4'b0010) begin
            S = 8'b01010111;
        end
    end
    if(A == 8'b01010110) begin
        if(B == 4'b0010) begin
            S = 8'b01011000;
        end
    end
    if(A == 8'b01010111) begin
        if(B == 4'b0010) begin
            S = 8'b01011001;
        end
    end
    if(A == 8'b01011000) begin
        if(B == 4'b0010) begin
            S = 8'b01011010;
        end
    end
    if(A == 8'b01011001) begin
        if(B == 4'b0010) begin
            S = 8'b01011011;
        end
    end
    if(A == 8'b01011010) begin
        if(B == 4'b0010) begin
            S = 8'b01011100;
        end
    end
    if(A == 8'b01011011) begin
        if(B == 4'b0010) begin
            S = 8'b01011101;
        end
    end
    if(A == 8'b01011100) begin
        if(B == 4'b0010) begin
            S = 8'b01011110;
        end
    end
    if(A == 8'b01011101) begin
        if(B == 4'b0010) begin
            S = 8'b01011111;
        end
    end
    if(A == 8'b01011110) begin
        if(B == 4'b0010) begin
            S = 8'b01100000;
        end
    end
    if(A == 8'b01011111) begin
        if(B == 4'b0010) begin
            S = 8'b01100001;
        end
    end
    if(A == 8'b01100000) begin
        if(B == 4'b0010) begin
            S = 8'b01100010;
        end
    end
    if(A == 8'b01100001) begin
        if(B == 4'b0010) begin
            S = 8'b01100011;
        end
    end
    if(A == 8'b00000000) begin
        if(B == 4'b0011) begin
            S = 8'b00000011;
        end
    end
    if(A == 8'b00000001) begin
        if(B == 4'b0011) begin
            S = 8'b00000100;
        end
    end
    if(A == 8'b00000010) begin
        if(B == 4'b0011) begin
            S = 8'b00000101;
        end
    end
    if(A == 8'b00000011) begin
        if(B == 4'b0011) begin
            S = 8'b00000110;
        end
    end
    if(A == 8'b00000100) begin
        if(B == 4'b0011) begin
            S = 8'b00000111;
        end
    end
    if(A == 8'b00000101) begin
        if(B == 4'b0011) begin
            S = 8'b00001000;
        end
    end
    if(A == 8'b00000110) begin
        if(B == 4'b0011) begin
            S = 8'b00001001;
        end
    end
    if(A == 8'b00000111) begin
        if(B == 4'b0011) begin
            S = 8'b00001010;
        end
    end
    if(A == 8'b00001000) begin
        if(B == 4'b0011) begin
            S = 8'b00001011;
        end
    end
    if(A == 8'b00001001) begin
        if(B == 4'b0011) begin
            S = 8'b00001100;
        end
    end
    if(A == 8'b00001010) begin
        if(B == 4'b0011) begin
            S = 8'b00001101;
        end
    end
    if(A == 8'b00001011) begin
        if(B == 4'b0011) begin
            S = 8'b00001110;
        end
    end
    if(A == 8'b00001100) begin
        if(B == 4'b0011) begin
            S = 8'b00001111;
        end
    end
    if(A == 8'b00001101) begin
        if(B == 4'b0011) begin
            S = 8'b00010000;
        end
    end
    if(A == 8'b00001110) begin
        if(B == 4'b0011) begin
            S = 8'b000010001;
        end
    end
    if(A == 8'b00001111) begin
        if(B == 4'b0011) begin
            S = 8'b000010010;
        end
    end
    if(A == 8'b00010000) begin
        if(B == 4'b0011) begin
            S = 8'b000010011;
        end
    end
    if(A == 8'b000010001) begin
        if(B == 4'b0011) begin
            S = 8'b000010100;
        end
    end
    if(A == 8'b000010010) begin
        if(B == 4'b0011) begin
            S = 8'b000010101;
        end
    end
    if(A == 8'b000010011) begin
        if(B == 4'b0011) begin
            S = 8'b000010110;
        end
    end
    if(A == 8'b000010100) begin
        if(B == 4'b0011) begin
            S = 8'b000010111;
        end
    end
    if(A == 8'b000010101) begin
        if(B == 4'b0011) begin
            S = 8'b00011000;
        end
    end
    if(A == 8'b000010110) begin
        if(B == 4'b0011) begin
            S = 8'b00011001;
        end
    end
    if(A == 8'b000010111) begin
        if(B == 4'b0011) begin
            S = 8'b00011010;
        end
    end
    if(A == 8'b00011000) begin
        if(B == 4'b0011) begin
            S = 8'b00011011;
        end
    end
    if(A == 8'b00011001) begin
        if(B == 4'b0011) begin
            S = 8'b00011100;
        end
    end
    if(A == 8'b00011010) begin
        if(B == 4'b0011) begin
            S = 8'b00011101;
        end
    end
    if(A == 8'b00011011) begin
        if(B == 4'b0011) begin
            S = 8'b00011110;
        end
    end
    if(A == 8'b00011100) begin
        if(B == 4'b0011) begin
            S = 8'b00011111;
        end
    end
    if(A == 8'b00011101) begin
        if(B == 4'b0011) begin
            S = 8'b00100000;
        end
    end
    if(A == 8'b00011110) begin
        if(B == 4'b0011) begin
            S = 8'b00100001;
        end
    end
    if(A == 8'b00011111) begin
        if(B == 4'b0011) begin
            S = 8'b00100010;
        end
    end
    if(A == 8'b00100000) begin
        if(B == 4'b0011) begin
            S = 8'b00100011;
        end
    end
    if(A == 8'b00100001) begin
        if(B == 4'b0011) begin
            S = 8'b00100100;
        end
    end
    if(A == 8'b00100010) begin
        if(B == 4'b0011) begin
            S = 8'b00100101;
        end
    end
    if(A == 8'b00100011) begin
        if(B == 4'b0011) begin
            S = 8'b00100110;
        end
    end
    if(A == 8'b00100100) begin
        if(B == 4'b0011) begin
            S = 8'b00100111;
        end
    end
    if(A == 8'b00100101) begin
        if(B == 4'b0011) begin
            S = 8'b00101000;
        end
    end
    if(A == 8'b00100110) begin
        if(B == 4'b0011) begin
            S = 8'b00101001;
        end
    end
    if(A == 8'b00100111) begin
        if(B == 4'b0011) begin
            S = 8'b00101010;
        end
    end
    if(A == 8'b00101000) begin
        if(B == 4'b0011) begin
            S = 8'b00101011;
        end
    end
    if(A == 8'b00101001) begin
        if(B == 4'b0011) begin
            S = 8'b00101100;
        end
    end
    if(A == 8'b00101010) begin
        if(B == 4'b0011) begin
            S = 8'b00101101;
        end
    end
    if(A == 8'b00101011) begin
        if(B == 4'b0011) begin
            S = 8'b00101110;
        end
    end
    if(A == 8'b00101100) begin
        if(B == 4'b0011) begin
            S = 8'b00101111;
        end
    end
    if(A == 8'b00101101) begin
        if(B == 4'b0011) begin
            S = 8'b00110000;
        end
    end
    if(A == 8'b00101110) begin
        if(B == 4'b0011) begin
            S = 8'b00110001;
        end
    end
    if(A == 8'b00101111) begin
        if(B == 4'b0011) begin
            S = 8'b00110010;
        end
    end
    if(A == 8'b00110000) begin
        if(B == 4'b0011) begin
            S = 8'b00110011;
        end
    end
    if(A == 8'b00110001) begin
        if(B == 4'b0011) begin
            S = 8'b00110100;
        end
    end
    if(A == 8'b00110010) begin
        if(B == 4'b0011) begin
            S = 8'b00110101;
        end
    end
    if(A == 8'b00110011) begin
        if(B == 4'b0011) begin
            S = 8'b00110110;
        end
    end
    if(A == 8'b00110100) begin
        if(B == 4'b0011) begin
            S = 8'b00110111;
        end
    end
    if(A == 8'b00110101) begin
        if(B == 4'b0011) begin
            S = 8'b00111000;
        end
    end
    if(A == 8'b00110110) begin
        if(B == 4'b0011) begin
            S = 8'b00111001;
        end
    end
    if(A == 8'b00110111) begin
        if(B == 4'b0011) begin
            S = 8'b00111010;
        end
    end
    if(A == 8'b00111000) begin
        if(B == 4'b0011) begin
            S = 8'b00111011;
        end
    end
    if(A == 8'b00111001) begin
        if(B == 4'b0011) begin
            S = 8'b00111100;
        end
    end
    if(A == 8'b00111010) begin
        if(B == 4'b0011) begin
            S = 8'b00111101;
        end
    end
    if(A == 8'b00111011) begin
        if(B == 4'b0011) begin
            S = 8'b00111110;
        end
    end
    if(A == 8'b00111100) begin
        if(B == 4'b0011) begin
            S = 8'b00111111;
        end
    end
    if(A == 8'b00111101) begin
        if(B == 4'b0011) begin
            S = 8'b01000000;
        end
    end
    if(A == 8'b00111110) begin
        if(B == 4'b0011) begin
            S = 8'b01000001;
        end
    end
    if(A == 8'b00111111) begin
        if(B == 4'b0011) begin
            S = 8'b01000010;
        end
    end
    if(A == 8'b01000000) begin
        if(B == 4'b0011) begin
            S = 8'b01000011;
        end
    end
    if(A == 8'b01000001) begin
        if(B == 4'b0011) begin
            S = 8'b01000100;
        end
    end
    if(A == 8'b01000010) begin
        if(B == 4'b0011) begin
            S = 8'b01000101;
        end
    end
    if(A == 8'b01000011) begin
        if(B == 4'b0011) begin
            S = 8'b01000110;
        end
    end
    if(A == 8'b01000100) begin
        if(B == 4'b0011) begin
            S = 8'b01000111;
        end
    end
    if(A == 8'b01000101) begin
        if(B == 4'b0011) begin
            S = 8'b01001000;
        end
    end
    if(A == 8'b01000110) begin
        if(B == 4'b0011) begin
            S = 8'b01001001;
        end
    end
    if(A == 8'b01000111) begin
        if(B == 4'b0011) begin
            S = 8'b01001010;
        end
    end
    if(A == 8'b01001000) begin
        if(B == 4'b0011) begin
            S = 8'b01001011;
        end
    end
    if(A == 8'b01001001) begin
        if(B == 4'b0011) begin
            S = 8'b01001100;
        end
    end
    if(A == 8'b01001010) begin
        if(B == 4'b0011) begin
            S = 8'b01001101;
        end
    end
    if(A == 8'b01001011) begin
        if(B == 4'b0011) begin
            S = 8'b01001110;
        end
    end
    if(A == 8'b01001100) begin
        if(B == 4'b0011) begin
            S = 8'b01001111;
        end
    end
    if(A == 8'b01001101) begin
        if(B == 4'b0011) begin
            S = 8'b01010000;
        end
    end
    if(A == 8'b01001110) begin
        if(B == 4'b0011) begin
            S = 8'b01010001;
        end
    end
    if(A == 8'b01001111) begin
        if(B == 4'b0011) begin
            S = 8'b01010010;
        end
    end
    if(A == 8'b01010000) begin
        if(B == 4'b0011) begin
            S = 8'b01010011;
        end
    end
    if(A == 8'b01010001) begin
        if(B == 4'b0011) begin
            S = 8'b01010100;
        end
    end
    if(A == 8'b01010010) begin
        if(B == 4'b0011) begin
            S = 8'b01010101;
        end
    end
    if(A == 8'b01010011) begin
        if(B == 4'b0011) begin
            S = 8'b01010110;
        end
    end
    if(A == 8'b01010100) begin
        if(B == 4'b0011) begin
            S = 8'b01010111;
        end
    end
    if(A == 8'b01010101) begin
        if(B == 4'b0011) begin
            S = 8'b01011000;
        end
    end
    if(A == 8'b01010110) begin
        if(B == 4'b0011) begin
            S = 8'b01011001;
        end
    end
    if(A == 8'b01010111) begin
        if(B == 4'b0011) begin
            S = 8'b01011010;
        end
    end
    if(A == 8'b01011000) begin
        if(B == 4'b0011) begin
            S = 8'b01011011;
        end
    end
    if(A == 8'b01011001) begin
        if(B == 4'b0011) begin
            S = 8'b01011100;
        end
    end
    if(A == 8'b01011010) begin
        if(B == 4'b0011) begin
            S = 8'b01011101;
        end
    end
    if(A == 8'b01011011) begin
        if(B == 4'b0011) begin
            S = 8'b01011110;
        end
    end
    if(A == 8'b01011100) begin
        if(B == 4'b0011) begin
            S = 8'b01011111;
        end
    end
    if(A == 8'b01011101) begin
        if(B == 4'b0011) begin
            S = 8'b01100000;
        end
    end
    if(A == 8'b01011110) begin
        if(B == 4'b0011) begin
            S = 8'b01100001;
        end
    end
    if(A == 8'b01011111) begin
        if(B == 4'b0011) begin
            S = 8'b01100010;
        end
    end
    if(A == 8'b01100000) begin
        if(B == 4'b0011) begin
            S = 8'b01100011;
        end
    end
    if(A == 8'b00000000) begin
        if(B == 4'b0100) begin
            S = 8'b00000100;
        end
    end
    if(A == 8'b00000001) begin
        if(B == 4'b0100) begin
            S = 8'b00000101;
        end
    end
    if(A == 8'b00000010) begin
        if(B == 4'b0100) begin
            S = 8'b00000110;
        end
    end
    if(A == 8'b00000011) begin
        if(B == 4'b0100) begin
            S = 8'b00000111;
        end
    end
    if(A == 8'b00000100) begin
        if(B == 4'b0100) begin
            S = 8'b00001000;
        end
    end
    if(A == 8'b00000101) begin
        if(B == 4'b0100) begin
            S = 8'b00001001;
        end
    end
    if(A == 8'b00000110) begin
        if(B == 4'b0100) begin
            S = 8'b00001010;
        end
    end
    if(A == 8'b00000111) begin
        if(B == 4'b0100) begin
            S = 8'b00001011;
        end
    end
    if(A == 8'b00001000) begin
        if(B == 4'b0100) begin
            S = 8'b00001100;
        end
    end
    if(A == 8'b00001001) begin
        if(B == 4'b0100) begin
            S = 8'b00001101;
        end
    end
    if(A == 8'b00001010) begin
        if(B == 4'b0100) begin
            S = 8'b00001110;
        end
    end
    if(A == 8'b00001011) begin
        if(B == 4'b0100) begin
            S = 8'b00001111;
        end
    end
    if(A == 8'b00001100) begin
        if(B == 4'b0100) begin
            S = 8'b00010000;
        end
    end
    if(A == 8'b00001101) begin
        if(B == 4'b0100) begin
            S = 8'b000010001;
        end
    end
    if(A == 8'b00001110) begin
        if(B == 4'b0100) begin
            S = 8'b000010010;
        end
    end
    if(A == 8'b00001111) begin
        if(B == 4'b0100) begin
            S = 8'b000010011;
        end
    end
    if(A == 8'b00010000) begin
        if(B == 4'b0100) begin
            S = 8'b000010100;
        end
    end
    if(A == 8'b000010001) begin
        if(B == 4'b0100) begin
            S = 8'b000010101;
        end
    end
    if(A == 8'b000010010) begin
        if(B == 4'b0100) begin
            S = 8'b000010110;
        end
    end
    if(A == 8'b000010011) begin
        if(B == 4'b0100) begin
            S = 8'b000010111;
        end
    end
    if(A == 8'b000010100) begin
        if(B == 4'b0100) begin
            S = 8'b00011000;
        end
    end
    if(A == 8'b000010101) begin
        if(B == 4'b0100) begin
            S = 8'b00011001;
        end
    end
    if(A == 8'b000010110) begin
        if(B == 4'b0100) begin
            S = 8'b00011010;
        end
    end
    if(A == 8'b000010111) begin
        if(B == 4'b0100) begin
            S = 8'b00011011;
        end
    end
    if(A == 8'b00011000) begin
        if(B == 4'b0100) begin
            S = 8'b00011100;
        end
    end
    if(A == 8'b00011001) begin
        if(B == 4'b0100) begin
            S = 8'b00011101;
        end
    end
    if(A == 8'b00011010) begin
        if(B == 4'b0100) begin
            S = 8'b00011110;
        end
    end
    if(A == 8'b00011011) begin
        if(B == 4'b0100) begin
            S = 8'b00011111;
        end
    end
    if(A == 8'b00011100) begin
        if(B == 4'b0100) begin
            S = 8'b00100000;
        end
    end
    if(A == 8'b00011101) begin
        if(B == 4'b0100) begin
            S = 8'b00100001;
        end
    end
    if(A == 8'b00011110) begin
        if(B == 4'b0100) begin
            S = 8'b00100010;
        end
    end
    if(A == 8'b00011111) begin
        if(B == 4'b0100) begin
            S = 8'b00100011;
        end
    end
    if(A == 8'b00100000) begin
        if(B == 4'b0100) begin
            S = 8'b00100100;
        end
    end
    if(A == 8'b00100001) begin
        if(B == 4'b0100) begin
            S = 8'b00100101;
        end
    end
    if(A == 8'b00100010) begin
        if(B == 4'b0100) begin
            S = 8'b00100110;
        end
    end
    if(A == 8'b00100011) begin
        if(B == 4'b0100) begin
            S = 8'b00100111;
        end
    end
    if(A == 8'b00100100) begin
        if(B == 4'b0100) begin
            S = 8'b00101000;
        end
    end
    if(A == 8'b00100101) begin
        if(B == 4'b0100) begin
            S = 8'b00101001;
        end
    end
    if(A == 8'b00100110) begin
        if(B == 4'b0100) begin
            S = 8'b00101010;
        end
    end
    if(A == 8'b00100111) begin
        if(B == 4'b0100) begin
            S = 8'b00101011;
        end
    end
    if(A == 8'b00101000) begin
        if(B == 4'b0100) begin
            S = 8'b00101100;
        end
    end
    if(A == 8'b00101001) begin
        if(B == 4'b0100) begin
            S = 8'b00101101;
        end
    end
    if(A == 8'b00101010) begin
        if(B == 4'b0100) begin
            S = 8'b00101110;
        end
    end
    if(A == 8'b00101011) begin
        if(B == 4'b0100) begin
            S = 8'b00101111;
        end
    end
    if(A == 8'b00101100) begin
        if(B == 4'b0100) begin
            S = 8'b00110000;
        end
    end
    if(A == 8'b00101101) begin
        if(B == 4'b0100) begin
            S = 8'b00110001;
        end
    end
    if(A == 8'b00101110) begin
        if(B == 4'b0100) begin
            S = 8'b00110010;
        end
    end
    if(A == 8'b00101111) begin
        if(B == 4'b0100) begin
            S = 8'b00110011;
        end
    end
    if(A == 8'b00110000) begin
        if(B == 4'b0100) begin
            S = 8'b00110100;
        end
    end
    if(A == 8'b00110001) begin
        if(B == 4'b0100) begin
            S = 8'b00110101;
        end
    end
    if(A == 8'b00110010) begin
        if(B == 4'b0100) begin
            S = 8'b00110110;
        end
    end
    if(A == 8'b00110011) begin
        if(B == 4'b0100) begin
            S = 8'b00110111;
        end
    end
    if(A == 8'b00110100) begin
        if(B == 4'b0100) begin
            S = 8'b00111000;
        end
    end
    if(A == 8'b00110101) begin
        if(B == 4'b0100) begin
            S = 8'b00111001;
        end
    end
    if(A == 8'b00110110) begin
        if(B == 4'b0100) begin
            S = 8'b00111010;
        end
    end
    if(A == 8'b00110111) begin
        if(B == 4'b0100) begin
            S = 8'b00111011;
        end
    end
    if(A == 8'b00111000) begin
        if(B == 4'b0100) begin
            S = 8'b00111100;
        end
    end
    if(A == 8'b00111001) begin
        if(B == 4'b0100) begin
            S = 8'b00111101;
        end
    end
    if(A == 8'b00111010) begin
        if(B == 4'b0100) begin
            S = 8'b00111110;
        end
    end
    if(A == 8'b00111011) begin
        if(B == 4'b0100) begin
            S = 8'b00111111;
        end
    end
    if(A == 8'b00111100) begin
        if(B == 4'b0100) begin
            S = 8'b01000000;
        end
    end
    if(A == 8'b00111101) begin
        if(B == 4'b0100) begin
            S = 8'b01000001;
        end
    end
    if(A == 8'b00111110) begin
        if(B == 4'b0100) begin
            S = 8'b01000010;
        end
    end
    if(A == 8'b00111111) begin
        if(B == 4'b0100) begin
            S = 8'b01000011;
        end
    end
    if(A == 8'b01000000) begin
        if(B == 4'b0100) begin
            S = 8'b01000100;
        end
    end
    if(A == 8'b01000001) begin
        if(B == 4'b0100) begin
            S = 8'b01000101;
        end
    end
    if(A == 8'b01000010) begin
        if(B == 4'b0100) begin
            S = 8'b01000110;
        end
    end
    if(A == 8'b01000011) begin
        if(B == 4'b0100) begin
            S = 8'b01000111;
        end
    end
    if(A == 8'b01000100) begin
        if(B == 4'b0100) begin
            S = 8'b01001000;
        end
    end
    if(A == 8'b01000101) begin
        if(B == 4'b0100) begin
            S = 8'b01001001;
        end
    end
    if(A == 8'b01000110) begin
        if(B == 4'b0100) begin
            S = 8'b01001010;
        end
    end
    if(A == 8'b01000111) begin
        if(B == 4'b0100) begin
            S = 8'b01001011;
        end
    end
    if(A == 8'b01001000) begin
        if(B == 4'b0100) begin
            S = 8'b01001100;
        end
    end
    if(A == 8'b01001001) begin
        if(B == 4'b0100) begin
            S = 8'b01001101;
        end
    end
    if(A == 8'b01001010) begin
        if(B == 4'b0100) begin
            S = 8'b01001110;
        end
    end
    if(A == 8'b01001011) begin
        if(B == 4'b0100) begin
            S = 8'b01001111;
        end
    end
    if(A == 8'b01001100) begin
        if(B == 4'b0100) begin
            S = 8'b01010000;
        end
    end
    if(A == 8'b01001101) begin
        if(B == 4'b0100) begin
            S = 8'b01010001;
        end
    end
    if(A == 8'b01001110) begin
        if(B == 4'b0100) begin
            S = 8'b01010010;
        end
    end
    if(A == 8'b01001111) begin
        if(B == 4'b0100) begin
            S = 8'b01010011;
        end
    end
    if(A == 8'b01010000) begin
        if(B == 4'b0100) begin
            S = 8'b01010100;
        end
    end
    if(A == 8'b01010001) begin
        if(B == 4'b0100) begin
            S = 8'b01010101;
        end
    end
    if(A == 8'b01010010) begin
        if(B == 4'b0100) begin
            S = 8'b01010110;
        end
    end
    if(A == 8'b01010011) begin
        if(B == 4'b0100) begin
            S = 8'b01010111;
        end
    end
    if(A == 8'b01010100) begin
        if(B == 4'b0100) begin
            S = 8'b01011000;
        end
    end
    if(A == 8'b01010101) begin
        if(B == 4'b0100) begin
            S = 8'b01011001;
        end
    end
    if(A == 8'b01010110) begin
        if(B == 4'b0100) begin
            S = 8'b01011010;
        end
    end
    if(A == 8'b01010111) begin
        if(B == 4'b0100) begin
            S = 8'b01011011;
        end
    end
    if(A == 8'b01011000) begin
        if(B == 4'b0100) begin
            S = 8'b01011100;
        end
    end
    if(A == 8'b01011001) begin
        if(B == 4'b0100) begin
            S = 8'b01011101;
        end
    end
    if(A == 8'b01011010) begin
        if(B == 4'b0100) begin
            S = 8'b01011110;
        end
    end
    if(A == 8'b01011011) begin
        if(B == 4'b0100) begin
            S = 8'b01011111;
        end
    end
    if(A == 8'b01011100) begin
        if(B == 4'b0100) begin
            S = 8'b01100000;
        end
    end
    if(A == 8'b01011101) begin
        if(B == 4'b0100) begin
            S = 8'b01100001;
        end
    end
    if(A == 8'b01011110) begin
        if(B == 4'b0100) begin
            S = 8'b01100010;
        end
    end
    if(A == 8'b01011111) begin
        if(B == 4'b0100) begin
            S = 8'b01100011;
        end
    end
    if(A == 8'b00000000) begin
        if(B == 4'b0101) begin
            S = 8'b00000101;
        end
    end
    if(A == 8'b00000001) begin
        if(B == 4'b0101) begin
            S = 8'b00000110;
        end
    end
    if(A == 8'b00000010) begin
        if(B == 4'b0101) begin
            S = 8'b00000111;
        end
    end
    if(A == 8'b00000011) begin
        if(B == 4'b0101) begin
            S = 8'b00001000;
        end
    end
    if(A == 8'b00000100) begin
        if(B == 4'b0101) begin
            S = 8'b00001001;
        end
    end
    if(A == 8'b00000101) begin
        if(B == 4'b0101) begin
            S = 8'b00001010;
        end
    end
    if(A == 8'b00000110) begin
        if(B == 4'b0101) begin
            S = 8'b00001011;
        end
    end
    if(A == 8'b00000111) begin
        if(B == 4'b0101) begin
            S = 8'b00001100;
        end
    end
    if(A == 8'b00001000) begin
        if(B == 4'b0101) begin
            S = 8'b00001101;
        end
    end
    if(A == 8'b00001001) begin
        if(B == 4'b0101) begin
            S = 8'b00001110;
        end
    end
    if(A == 8'b00001010) begin
        if(B == 4'b0101) begin
            S = 8'b00001111;
        end
    end
    if(A == 8'b00001011) begin
        if(B == 4'b0101) begin
            S = 8'b00010000;
        end
    end
    if(A == 8'b00001100) begin
        if(B == 4'b0101) begin
            S = 8'b000010001;
        end
    end
    if(A == 8'b00001101) begin
        if(B == 4'b0101) begin
            S = 8'b000010010;
        end
    end
    if(A == 8'b00001110) begin
        if(B == 4'b0101) begin
            S = 8'b000010011;
        end
    end
    if(A == 8'b00001111) begin
        if(B == 4'b0101) begin
            S = 8'b000010100;
        end
    end
    if(A == 8'b00010000) begin
        if(B == 4'b0101) begin
            S = 8'b000010101;
        end
    end
    if(A == 8'b000010001) begin
        if(B == 4'b0101) begin
            S = 8'b000010110;
        end
    end
    if(A == 8'b000010010) begin
        if(B == 4'b0101) begin
            S = 8'b000010111;
        end
    end
    if(A == 8'b000010011) begin
        if(B == 4'b0101) begin
            S = 8'b00011000;
        end
    end
    if(A == 8'b000010100) begin
        if(B == 4'b0101) begin
            S = 8'b00011001;
        end
    end
    if(A == 8'b000010101) begin
        if(B == 4'b0101) begin
            S = 8'b00011010;
        end
    end
    if(A == 8'b000010110) begin
        if(B == 4'b0101) begin
            S = 8'b00011011;
        end
    end
    if(A == 8'b000010111) begin
        if(B == 4'b0101) begin
            S = 8'b00011100;
        end
    end
    if(A == 8'b00011000) begin
        if(B == 4'b0101) begin
            S = 8'b00011101;
        end
    end
    if(A == 8'b00011001) begin
        if(B == 4'b0101) begin
            S = 8'b00011110;
        end
    end
    if(A == 8'b00011010) begin
        if(B == 4'b0101) begin
            S = 8'b00011111;
        end
    end
    if(A == 8'b00011011) begin
        if(B == 4'b0101) begin
            S = 8'b00100000;
        end
    end
    if(A == 8'b00011100) begin
        if(B == 4'b0101) begin
            S = 8'b00100001;
        end
    end
    if(A == 8'b00011101) begin
        if(B == 4'b0101) begin
            S = 8'b00100010;
        end
    end
    if(A == 8'b00011110) begin
        if(B == 4'b0101) begin
            S = 8'b00100011;
        end
    end
    if(A == 8'b00011111) begin
        if(B == 4'b0101) begin
            S = 8'b00100100;
        end
    end
    if(A == 8'b00100000) begin
        if(B == 4'b0101) begin
            S = 8'b00100101;
        end
    end
    if(A == 8'b00100001) begin
        if(B == 4'b0101) begin
            S = 8'b00100110;
        end
    end
    if(A == 8'b00100010) begin
        if(B == 4'b0101) begin
            S = 8'b00100111;
        end
    end
    if(A == 8'b00100011) begin
        if(B == 4'b0101) begin
            S = 8'b00101000;
        end
    end
    if(A == 8'b00100100) begin
        if(B == 4'b0101) begin
            S = 8'b00101001;
        end
    end
    if(A == 8'b00100101) begin
        if(B == 4'b0101) begin
            S = 8'b00101010;
        end
    end
    if(A == 8'b00100110) begin
        if(B == 4'b0101) begin
            S = 8'b00101011;
        end
    end
    if(A == 8'b00100111) begin
        if(B == 4'b0101) begin
            S = 8'b00101100;
        end
    end
    if(A == 8'b00101000) begin
        if(B == 4'b0101) begin
            S = 8'b00101101;
        end
    end
    if(A == 8'b00101001) begin
        if(B == 4'b0101) begin
            S = 8'b00101110;
        end
    end
    if(A == 8'b00101010) begin
        if(B == 4'b0101) begin
            S = 8'b00101111;
        end
    end
    if(A == 8'b00101011) begin
        if(B == 4'b0101) begin
            S = 8'b00110000;
        end
    end
    if(A == 8'b00101100) begin
        if(B == 4'b0101) begin
            S = 8'b00110001;
        end
    end
    if(A == 8'b00101101) begin
        if(B == 4'b0101) begin
            S = 8'b00110010;
        end
    end
    if(A == 8'b00101110) begin
        if(B == 4'b0101) begin
            S = 8'b00110011;
        end
    end
    if(A == 8'b00101111) begin
        if(B == 4'b0101) begin
            S = 8'b00110100;
        end
    end
    if(A == 8'b00110000) begin
        if(B == 4'b0101) begin
            S = 8'b00110101;
        end
    end
    if(A == 8'b00110001) begin
        if(B == 4'b0101) begin
            S = 8'b00110110;
        end
    end
    if(A == 8'b00110010) begin
        if(B == 4'b0101) begin
            S = 8'b00110111;
        end
    end
    if(A == 8'b00110011) begin
        if(B == 4'b0101) begin
            S = 8'b00111000;
        end
    end
    if(A == 8'b00110100) begin
        if(B == 4'b0101) begin
            S = 8'b00111001;
        end
    end
    if(A == 8'b00110101) begin
        if(B == 4'b0101) begin
            S = 8'b00111010;
        end
    end
    if(A == 8'b00110110) begin
        if(B == 4'b0101) begin
            S = 8'b00111011;
        end
    end
    if(A == 8'b00110111) begin
        if(B == 4'b0101) begin
            S = 8'b00111100;
        end
    end
    if(A == 8'b00111000) begin
        if(B == 4'b0101) begin
            S = 8'b00111101;
        end
    end
    if(A == 8'b00111001) begin
        if(B == 4'b0101) begin
            S = 8'b00111110;
        end
    end
    if(A == 8'b00111010) begin
        if(B == 4'b0101) begin
            S = 8'b00111111;
        end
    end
    if(A == 8'b00111011) begin
        if(B == 4'b0101) begin
            S = 8'b01000000;
        end
    end
    if(A == 8'b00111100) begin
        if(B == 4'b0101) begin
            S = 8'b01000001;
        end
    end
    if(A == 8'b00111101) begin
        if(B == 4'b0101) begin
            S = 8'b01000010;
        end
    end
    if(A == 8'b00111110) begin
        if(B == 4'b0101) begin
            S = 8'b01000011;
        end
    end
    if(A == 8'b00111111) begin
        if(B == 4'b0101) begin
            S = 8'b01000100;
        end
    end
    if(A == 8'b01000000) begin
        if(B == 4'b0101) begin
            S = 8'b01000101;
        end
    end
    if(A == 8'b01000001) begin
        if(B == 4'b0101) begin
            S = 8'b01000110;
        end
    end
    if(A == 8'b01000010) begin
        if(B == 4'b0101) begin
            S = 8'b01000111;
        end
    end
    if(A == 8'b01000011) begin
        if(B == 4'b0101) begin
            S = 8'b01001000;
        end
    end
    if(A == 8'b01000100) begin
        if(B == 4'b0101) begin
            S = 8'b01001001;
        end
    end
    if(A == 8'b01000101) begin
        if(B == 4'b0101) begin
            S = 8'b01001010;
        end
    end
    if(A == 8'b01000110) begin
        if(B == 4'b0101) begin
            S = 8'b01001011;
        end
    end
    if(A == 8'b01000111) begin
        if(B == 4'b0101) begin
            S = 8'b01001100;
        end
    end
    if(A == 8'b01001000) begin
        if(B == 4'b0101) begin
            S = 8'b01001101;
        end
    end
    if(A == 8'b01001001) begin
        if(B == 4'b0101) begin
            S = 8'b01001110;
        end
    end
    if(A == 8'b01001010) begin
        if(B == 4'b0101) begin
            S = 8'b01001111;
        end
    end
    if(A == 8'b01001011) begin
        if(B == 4'b0101) begin
            S = 8'b01010000;
        end
    end
    if(A == 8'b01001100) begin
        if(B == 4'b0101) begin
            S = 8'b01010001;
        end
    end
    if(A == 8'b01001101) begin
        if(B == 4'b0101) begin
            S = 8'b01010010;
        end
    end
    if(A == 8'b01001110) begin
        if(B == 4'b0101) begin
            S = 8'b01010011;
        end
    end
    if(A == 8'b01001111) begin
        if(B == 4'b0101) begin
            S = 8'b01010100;
        end
    end
    if(A == 8'b01010000) begin
        if(B == 4'b0101) begin
            S = 8'b01010101;
        end
    end
    if(A == 8'b01010001) begin
        if(B == 4'b0101) begin
            S = 8'b01010110;
        end
    end
    if(A == 8'b01010010) begin
        if(B == 4'b0101) begin
            S = 8'b01010111;
        end
    end
    if(A == 8'b01010011) begin
        if(B == 4'b0101) begin
            S = 8'b01011000;
        end
    end
    if(A == 8'b01010100) begin
        if(B == 4'b0101) begin
            S = 8'b01011001;
        end
    end
    if(A == 8'b01010101) begin
        if(B == 4'b0101) begin
            S = 8'b01011010;
        end
    end
    if(A == 8'b01010110) begin
        if(B == 4'b0101) begin
            S = 8'b01011011;
        end
    end
    if(A == 8'b01010111) begin
        if(B == 4'b0101) begin
            S = 8'b01011100;
        end
    end
    if(A == 8'b01011000) begin
        if(B == 4'b0101) begin
            S = 8'b01011101;
        end
    end
    if(A == 8'b01011001) begin
        if(B == 4'b0101) begin
            S = 8'b01011110;
        end
    end
    if(A == 8'b01011010) begin
        if(B == 4'b0101) begin
            S = 8'b01011111;
        end
    end
    if(A == 8'b01011011) begin
        if(B == 4'b0101) begin
            S = 8'b01100000;
        end
    end
    if(A == 8'b01011100) begin
        if(B == 4'b0101) begin
            S = 8'b01100001;
        end
    end
    if(A == 8'b01011101) begin
        if(B == 4'b0101) begin
            S = 8'b01100010;
        end
    end
    if(A == 8'b01011110) begin
        if(B == 4'b0101) begin
            S = 8'b01100011;
        end
    end
    if(A == 8'b00000000) begin
        if(B == 4'b0110) begin
            S = 8'b00000110;
        end
    end
    if(A == 8'b00000001) begin
        if(B == 4'b0110) begin
            S = 8'b00000111;
        end
    end
    if(A == 8'b00000010) begin
        if(B == 4'b0110) begin
            S = 8'b00001000;
        end
    end
    if(A == 8'b00000011) begin
        if(B == 4'b0110) begin
            S = 8'b00001001;
        end
    end
    if(A == 8'b00000100) begin
        if(B == 4'b0110) begin
            S = 8'b00001010;
        end
    end
    if(A == 8'b00000101) begin
        if(B == 4'b0110) begin
            S = 8'b00001011;
        end
    end
    if(A == 8'b00000110) begin
        if(B == 4'b0110) begin
            S = 8'b00001100;
        end
    end
    if(A == 8'b00000111) begin
        if(B == 4'b0110) begin
            S = 8'b00001101;
        end
    end
    if(A == 8'b00001000) begin
        if(B == 4'b0110) begin
            S = 8'b00001110;
        end
    end
    if(A == 8'b00001001) begin
        if(B == 4'b0110) begin
            S = 8'b00001111;
        end
    end
    if(A == 8'b00001010) begin
        if(B == 4'b0110) begin
            S = 8'b00010000;
        end
    end
    if(A == 8'b00001011) begin
        if(B == 4'b0110) begin
            S = 8'b000010001;
        end
    end
    if(A == 8'b00001100) begin
        if(B == 4'b0110) begin
            S = 8'b000010010;
        end
    end
    if(A == 8'b00001101) begin
        if(B == 4'b0110) begin
            S = 8'b000010011;
        end
    end
    if(A == 8'b00001110) begin
        if(B == 4'b0110) begin
            S = 8'b000010100;
        end
    end
    if(A == 8'b00001111) begin
        if(B == 4'b0110) begin
            S = 8'b000010101;
        end
    end
    if(A == 8'b00010000) begin
        if(B == 4'b0110) begin
            S = 8'b000010110;
        end
    end
    if(A == 8'b000010001) begin
        if(B == 4'b0110) begin
            S = 8'b000010111;
        end
    end
    if(A == 8'b000010010) begin
        if(B == 4'b0110) begin
            S = 8'b00011000;
        end
    end
    if(A == 8'b000010011) begin
        if(B == 4'b0110) begin
            S = 8'b00011001;
        end
    end
    if(A == 8'b000010100) begin
        if(B == 4'b0110) begin
            S = 8'b00011010;
        end
    end
    if(A == 8'b000010101) begin
        if(B == 4'b0110) begin
            S = 8'b00011011;
        end
    end
    if(A == 8'b000010110) begin
        if(B == 4'b0110) begin
            S = 8'b00011100;
        end
    end
    if(A == 8'b000010111) begin
        if(B == 4'b0110) begin
            S = 8'b00011101;
        end
    end
    if(A == 8'b00011000) begin
        if(B == 4'b0110) begin
            S = 8'b00011110;
        end
    end
    if(A == 8'b00011001) begin
        if(B == 4'b0110) begin
            S = 8'b00011111;
        end
    end
    if(A == 8'b00011010) begin
        if(B == 4'b0110) begin
            S = 8'b00100000;
        end
    end
    if(A == 8'b00011011) begin
        if(B == 4'b0110) begin
            S = 8'b00100001;
        end
    end
    if(A == 8'b00011100) begin
        if(B == 4'b0110) begin
            S = 8'b00100010;
        end
    end
    if(A == 8'b00011101) begin
        if(B == 4'b0110) begin
            S = 8'b00100011;
        end
    end
    if(A == 8'b00011110) begin
        if(B == 4'b0110) begin
            S = 8'b00100100;
        end
    end
    if(A == 8'b00011111) begin
        if(B == 4'b0110) begin
            S = 8'b00100101;
        end
    end
    if(A == 8'b00100000) begin
        if(B == 4'b0110) begin
            S = 8'b00100110;
        end
    end
    if(A == 8'b00100001) begin
        if(B == 4'b0110) begin
            S = 8'b00100111;
        end
    end
    if(A == 8'b00100010) begin
        if(B == 4'b0110) begin
            S = 8'b00101000;
        end
    end
    if(A == 8'b00100011) begin
        if(B == 4'b0110) begin
            S = 8'b00101001;
        end
    end
    if(A == 8'b00100100) begin
        if(B == 4'b0110) begin
            S = 8'b00101010;
        end
    end
    if(A == 8'b00100101) begin
        if(B == 4'b0110) begin
            S = 8'b00101011;
        end
    end
    if(A == 8'b00100110) begin
        if(B == 4'b0110) begin
            S = 8'b00101100;
        end
    end
    if(A == 8'b00100111) begin
        if(B == 4'b0110) begin
            S = 8'b00101101;
        end
    end
    if(A == 8'b00101000) begin
        if(B == 4'b0110) begin
            S = 8'b00101110;
        end
    end
    if(A == 8'b00101001) begin
        if(B == 4'b0110) begin
            S = 8'b00101111;
        end
    end
    if(A == 8'b00101010) begin
        if(B == 4'b0110) begin
            S = 8'b00110000;
        end
    end
    if(A == 8'b00101011) begin
        if(B == 4'b0110) begin
            S = 8'b00110001;
        end
    end
    if(A == 8'b00101100) begin
        if(B == 4'b0110) begin
            S = 8'b00110010;
        end
    end
    if(A == 8'b00101101) begin
        if(B == 4'b0110) begin
            S = 8'b00110011;
        end
    end
    if(A == 8'b00101110) begin
        if(B == 4'b0110) begin
            S = 8'b00110100;
        end
    end
    if(A == 8'b00101111) begin
        if(B == 4'b0110) begin
            S = 8'b00110101;
        end
    end
    if(A == 8'b00110000) begin
        if(B == 4'b0110) begin
            S = 8'b00110110;
        end
    end
    if(A == 8'b00110001) begin
        if(B == 4'b0110) begin
            S = 8'b00110111;
        end
    end
    if(A == 8'b00110010) begin
        if(B == 4'b0110) begin
            S = 8'b00111000;
        end
    end
    if(A == 8'b00110011) begin
        if(B == 4'b0110) begin
            S = 8'b00111001;
        end
    end
    if(A == 8'b00110100) begin
        if(B == 4'b0110) begin
            S = 8'b00111010;
        end
    end
    if(A == 8'b00110101) begin
        if(B == 4'b0110) begin
            S = 8'b00111011;
        end
    end
    if(A == 8'b00110110) begin
        if(B == 4'b0110) begin
            S = 8'b00111100;
        end
    end
    if(A == 8'b00110111) begin
        if(B == 4'b0110) begin
            S = 8'b00111101;
        end
    end
    if(A == 8'b00111000) begin
        if(B == 4'b0110) begin
            S = 8'b00111110;
        end
    end
    if(A == 8'b00111001) begin
        if(B == 4'b0110) begin
            S = 8'b00111111;
        end
    end
    if(A == 8'b00111010) begin
        if(B == 4'b0110) begin
            S = 8'b01000000;
        end
    end
    if(A == 8'b00111011) begin
        if(B == 4'b0110) begin
            S = 8'b01000001;
        end
    end
    if(A == 8'b00111100) begin
        if(B == 4'b0110) begin
            S = 8'b01000010;
        end
    end
    if(A == 8'b00111101) begin
        if(B == 4'b0110) begin
            S = 8'b01000011;
        end
    end
    if(A == 8'b00111110) begin
        if(B == 4'b0110) begin
            S = 8'b01000100;
        end
    end
    if(A == 8'b00111111) begin
        if(B == 4'b0110) begin
            S = 8'b01000101;
        end
    end
    if(A == 8'b01000000) begin
        if(B == 4'b0110) begin
            S = 8'b01000110;
        end
    end
    if(A == 8'b01000001) begin
        if(B == 4'b0110) begin
            S = 8'b01000111;
        end
    end
    if(A == 8'b01000010) begin
        if(B == 4'b0110) begin
            S = 8'b01001000;
        end
    end
    if(A == 8'b01000011) begin
        if(B == 4'b0110) begin
            S = 8'b01001001;
        end
    end
    if(A == 8'b01000100) begin
        if(B == 4'b0110) begin
            S = 8'b01001010;
        end
    end
    if(A == 8'b01000101) begin
        if(B == 4'b0110) begin
            S = 8'b01001011;
        end
    end
    if(A == 8'b01000110) begin
        if(B == 4'b0110) begin
            S = 8'b01001100;
        end
    end
    if(A == 8'b01000111) begin
        if(B == 4'b0110) begin
            S = 8'b01001101;
        end
    end
    if(A == 8'b01001000) begin
        if(B == 4'b0110) begin
            S = 8'b01001110;
        end
    end
    if(A == 8'b01001001) begin
        if(B == 4'b0110) begin
            S = 8'b01001111;
        end
    end
    if(A == 8'b01001010) begin
        if(B == 4'b0110) begin
            S = 8'b01010000;
        end
    end
    if(A == 8'b01001011) begin
        if(B == 4'b0110) begin
            S = 8'b01010001;
        end
    end
    if(A == 8'b01001100) begin
        if(B == 4'b0110) begin
            S = 8'b01010010;
        end
    end
    if(A == 8'b01001101) begin
        if(B == 4'b0110) begin
            S = 8'b01010011;
        end
    end
    if(A == 8'b01001110) begin
        if(B == 4'b0110) begin
            S = 8'b01010100;
        end
    end
    if(A == 8'b01001111) begin
        if(B == 4'b0110) begin
            S = 8'b01010101;
        end
    end
    if(A == 8'b01010000) begin
        if(B == 4'b0110) begin
            S = 8'b01010110;
        end
    end
    if(A == 8'b01010001) begin
        if(B == 4'b0110) begin
            S = 8'b01010111;
        end
    end
    if(A == 8'b01010010) begin
        if(B == 4'b0110) begin
            S = 8'b01011000;
        end
    end
    if(A == 8'b01010011) begin
        if(B == 4'b0110) begin
            S = 8'b01011001;
        end
    end
    if(A == 8'b01010100) begin
        if(B == 4'b0110) begin
            S = 8'b01011010;
        end
    end
    if(A == 8'b01010101) begin
        if(B == 4'b0110) begin
            S = 8'b01011011;
        end
    end
    if(A == 8'b01010110) begin
        if(B == 4'b0110) begin
            S = 8'b01011100;
        end
    end
    if(A == 8'b01010111) begin
        if(B == 4'b0110) begin
            S = 8'b01011101;
        end
    end
    if(A == 8'b01011000) begin
        if(B == 4'b0110) begin
            S = 8'b01011110;
        end
    end
    if(A == 8'b01011001) begin
        if(B == 4'b0110) begin
            S = 8'b01011111;
        end
    end
    if(A == 8'b01011010) begin
        if(B == 4'b0110) begin
            S = 8'b01100000;
        end
    end
    if(A == 8'b01011011) begin
        if(B == 4'b0110) begin
            S = 8'b01100001;
        end
    end
    if(A == 8'b01011100) begin
        if(B == 4'b0110) begin
            S = 8'b01100010;
        end
    end
    if(A == 8'b01011101) begin
        if(B == 4'b0110) begin
            S = 8'b01100011;
        end
    end
    if(A == 8'b00000000) begin
        if(B == 4'b0111) begin
            S = 8'b00000111;
        end
    end
    if(A == 8'b00000001) begin
        if(B == 4'b0111) begin
            S = 8'b00001000;
        end
    end
    if(A == 8'b00000010) begin
        if(B == 4'b0111) begin
            S = 8'b00001001;
        end
    end
    if(A == 8'b00000011) begin
        if(B == 4'b0111) begin
            S = 8'b00001010;
        end
    end
    if(A == 8'b00000100) begin
        if(B == 4'b0111) begin
            S = 8'b00001011;
        end
    end
    if(A == 8'b00000101) begin
        if(B == 4'b0111) begin
            S = 8'b00001100;
        end
    end
    if(A == 8'b00000110) begin
        if(B == 4'b0111) begin
            S = 8'b00001101;
        end
    end
    if(A == 8'b00000111) begin
        if(B == 4'b0111) begin
            S = 8'b00001110;
        end
    end
    if(A == 8'b00001000) begin
        if(B == 4'b0111) begin
            S = 8'b00001111;
        end
    end
    if(A == 8'b00001001) begin
        if(B == 4'b0111) begin
            S = 8'b00010000;
        end
    end
    if(A == 8'b00001010) begin
        if(B == 4'b0111) begin
            S = 8'b000010001;
        end
    end
    if(A == 8'b00001011) begin
        if(B == 4'b0111) begin
            S = 8'b000010010;
        end
    end
    if(A == 8'b00001100) begin
        if(B == 4'b0111) begin
            S = 8'b000010011;
        end
    end
    if(A == 8'b00001101) begin
        if(B == 4'b0111) begin
            S = 8'b000010100;
        end
    end
    if(A == 8'b00001110) begin
        if(B == 4'b0111) begin
            S = 8'b000010101;
        end
    end
    if(A == 8'b00001111) begin
        if(B == 4'b0111) begin
            S = 8'b000010110;
        end
    end
    if(A == 8'b00010000) begin
        if(B == 4'b0111) begin
            S = 8'b000010111;
        end
    end
    if(A == 8'b000010001) begin
        if(B == 4'b0111) begin
            S = 8'b00011000;
        end
    end
    if(A == 8'b000010010) begin
        if(B == 4'b0111) begin
            S = 8'b00011001;
        end
    end
    if(A == 8'b000010011) begin
        if(B == 4'b0111) begin
            S = 8'b00011010;
        end
    end
    if(A == 8'b000010100) begin
        if(B == 4'b0111) begin
            S = 8'b00011011;
        end
    end
    if(A == 8'b000010101) begin
        if(B == 4'b0111) begin
            S = 8'b00011100;
        end
    end
    if(A == 8'b000010110) begin
        if(B == 4'b0111) begin
            S = 8'b00011101;
        end
    end
    if(A == 8'b000010111) begin
        if(B == 4'b0111) begin
            S = 8'b00011110;
        end
    end
    if(A == 8'b00011000) begin
        if(B == 4'b0111) begin
            S = 8'b00011111;
        end
    end
    if(A == 8'b00011001) begin
        if(B == 4'b0111) begin
            S = 8'b00100000;
        end
    end
    if(A == 8'b00011010) begin
        if(B == 4'b0111) begin
            S = 8'b00100001;
        end
    end
    if(A == 8'b00011011) begin
        if(B == 4'b0111) begin
            S = 8'b00100010;
        end
    end
    if(A == 8'b00011100) begin
        if(B == 4'b0111) begin
            S = 8'b00100011;
        end
    end
    if(A == 8'b00011101) begin
        if(B == 4'b0111) begin
            S = 8'b00100100;
        end
    end
    if(A == 8'b00011110) begin
        if(B == 4'b0111) begin
            S = 8'b00100101;
        end
    end
    if(A == 8'b00011111) begin
        if(B == 4'b0111) begin
            S = 8'b00100110;
        end
    end
    if(A == 8'b00100000) begin
        if(B == 4'b0111) begin
            S = 8'b00100111;
        end
    end
    if(A == 8'b00100001) begin
        if(B == 4'b0111) begin
            S = 8'b00101000;
        end
    end
    if(A == 8'b00100010) begin
        if(B == 4'b0111) begin
            S = 8'b00101001;
        end
    end
    if(A == 8'b00100011) begin
        if(B == 4'b0111) begin
            S = 8'b00101010;
        end
    end
    if(A == 8'b00100100) begin
        if(B == 4'b0111) begin
            S = 8'b00101011;
        end
    end
    if(A == 8'b00100101) begin
        if(B == 4'b0111) begin
            S = 8'b00101100;
        end
    end
    if(A == 8'b00100110) begin
        if(B == 4'b0111) begin
            S = 8'b00101101;
        end
    end
    if(A == 8'b00100111) begin
        if(B == 4'b0111) begin
            S = 8'b00101110;
        end
    end
    if(A == 8'b00101000) begin
        if(B == 4'b0111) begin
            S = 8'b00101111;
        end
    end
    if(A == 8'b00101001) begin
        if(B == 4'b0111) begin
            S = 8'b00110000;
        end
    end
    if(A == 8'b00101010) begin
        if(B == 4'b0111) begin
            S = 8'b00110001;
        end
    end
    if(A == 8'b00101011) begin
        if(B == 4'b0111) begin
            S = 8'b00110010;
        end
    end
    if(A == 8'b00101100) begin
        if(B == 4'b0111) begin
            S = 8'b00110011;
        end
    end
    if(A == 8'b00101101) begin
        if(B == 4'b0111) begin
            S = 8'b00110100;
        end
    end
    if(A == 8'b00101110) begin
        if(B == 4'b0111) begin
            S = 8'b00110101;
        end
    end
    if(A == 8'b00101111) begin
        if(B == 4'b0111) begin
            S = 8'b00110110;
        end
    end
    if(A == 8'b00110000) begin
        if(B == 4'b0111) begin
            S = 8'b00110111;
        end
    end
    if(A == 8'b00110001) begin
        if(B == 4'b0111) begin
            S = 8'b00111000;
        end
    end
    if(A == 8'b00110010) begin
        if(B == 4'b0111) begin
            S = 8'b00111001;
        end
    end
    if(A == 8'b00110011) begin
        if(B == 4'b0111) begin
            S = 8'b00111010;
        end
    end
    if(A == 8'b00110100) begin
        if(B == 4'b0111) begin
            S = 8'b00111011;
        end
    end
    if(A == 8'b00110101) begin
        if(B == 4'b0111) begin
            S = 8'b00111100;
        end
    end
    if(A == 8'b00110110) begin
        if(B == 4'b0111) begin
            S = 8'b00111101;
        end
    end
    if(A == 8'b00110111) begin
        if(B == 4'b0111) begin
            S = 8'b00111110;
        end
    end
    if(A == 8'b00111000) begin
        if(B == 4'b0111) begin
            S = 8'b00111111;
        end
    end
    if(A == 8'b00111001) begin
        if(B == 4'b0111) begin
            S = 8'b01000000;
        end
    end
    if(A == 8'b00111010) begin
        if(B == 4'b0111) begin
            S = 8'b01000001;
        end
    end
    if(A == 8'b00111011) begin
        if(B == 4'b0111) begin
            S = 8'b01000010;
        end
    end
    if(A == 8'b00111100) begin
        if(B == 4'b0111) begin
            S = 8'b01000011;
        end
    end
    if(A == 8'b00111101) begin
        if(B == 4'b0111) begin
            S = 8'b01000100;
        end
    end
    if(A == 8'b00111110) begin
        if(B == 4'b0111) begin
            S = 8'b01000101;
        end
    end
    if(A == 8'b00111111) begin
        if(B == 4'b0111) begin
            S = 8'b01000110;
        end
    end
    if(A == 8'b01000000) begin
        if(B == 4'b0111) begin
            S = 8'b01000111;
        end
    end
    if(A == 8'b01000001) begin
        if(B == 4'b0111) begin
            S = 8'b01001000;
        end
    end
    if(A == 8'b01000010) begin
        if(B == 4'b0111) begin
            S = 8'b01001001;
        end
    end
    if(A == 8'b01000011) begin
        if(B == 4'b0111) begin
            S = 8'b01001010;
        end
    end
    if(A == 8'b01000100) begin
        if(B == 4'b0111) begin
            S = 8'b01001011;
        end
    end
    if(A == 8'b01000101) begin
        if(B == 4'b0111) begin
            S = 8'b01001100;
        end
    end
    if(A == 8'b01000110) begin
        if(B == 4'b0111) begin
            S = 8'b01001101;
        end
    end
    if(A == 8'b01000111) begin
        if(B == 4'b0111) begin
            S = 8'b01001110;
        end
    end
    if(A == 8'b01001000) begin
        if(B == 4'b0111) begin
            S = 8'b01001111;
        end
    end
    if(A == 8'b01001001) begin
        if(B == 4'b0111) begin
            S = 8'b01010000;
        end
    end
    if(A == 8'b01001010) begin
        if(B == 4'b0111) begin
            S = 8'b01010001;
        end
    end
    if(A == 8'b01001011) begin
        if(B == 4'b0111) begin
            S = 8'b01010010;
        end
    end
    if(A == 8'b01001100) begin
        if(B == 4'b0111) begin
            S = 8'b01010011;
        end
    end
    if(A == 8'b01001101) begin
        if(B == 4'b0111) begin
            S = 8'b01010100;
        end
    end
    if(A == 8'b01001110) begin
        if(B == 4'b0111) begin
            S = 8'b01010101;
        end
    end
    if(A == 8'b01001111) begin
        if(B == 4'b0111) begin
            S = 8'b01010110;
        end
    end
    if(A == 8'b01010000) begin
        if(B == 4'b0111) begin
            S = 8'b01010111;
        end
    end
    if(A == 8'b01010001) begin
        if(B == 4'b0111) begin
            S = 8'b01011000;
        end
    end
    if(A == 8'b01010010) begin
        if(B == 4'b0111) begin
            S = 8'b01011001;
        end
    end
    if(A == 8'b01010011) begin
        if(B == 4'b0111) begin
            S = 8'b01011010;
        end
    end
    if(A == 8'b01010100) begin
        if(B == 4'b0111) begin
            S = 8'b01011011;
        end
    end
    if(A == 8'b01010101) begin
        if(B == 4'b0111) begin
            S = 8'b01011100;
        end
    end
    if(A == 8'b01010110) begin
        if(B == 4'b0111) begin
            S = 8'b01011101;
        end
    end
    if(A == 8'b01010111) begin
        if(B == 4'b0111) begin
            S = 8'b01011110;
        end
    end
    if(A == 8'b01011000) begin
        if(B == 4'b0111) begin
            S = 8'b01011111;
        end
    end
    if(A == 8'b01011001) begin
        if(B == 4'b0111) begin
            S = 8'b01100000;
        end
    end
    if(A == 8'b01011010) begin
        if(B == 4'b0111) begin
            S = 8'b01100001;
        end
    end
    if(A == 8'b01011011) begin
        if(B == 4'b0111) begin
            S = 8'b01100010;
        end
    end
    if(A == 8'b01011100) begin
        if(B == 4'b0111) begin
            S = 8'b01100011;
        end
    end
    if(A == 8'b00000000) begin
        if(B == 4'b1000) begin
            S = 8'b00001000;
        end
    end
    if(A == 8'b00000001) begin
        if(B == 4'b1000) begin
            S = 8'b00001001;
        end
    end
    if(A == 8'b00000010) begin
        if(B == 4'b1000) begin
            S = 8'b00001010;
        end
    end
    if(A == 8'b00000011) begin
        if(B == 4'b1000) begin
            S = 8'b00001011;
        end
    end
    if(A == 8'b00000100) begin
        if(B == 4'b1000) begin
            S = 8'b00001100;
        end
    end
    if(A == 8'b00000101) begin
        if(B == 4'b1000) begin
            S = 8'b00001101;
        end
    end
    if(A == 8'b00000110) begin
        if(B == 4'b1000) begin
            S = 8'b00001110;
        end
    end
    if(A == 8'b00000111) begin
        if(B == 4'b1000) begin
            S = 8'b00001111;
        end
    end
    if(A == 8'b00001000) begin
        if(B == 4'b1000) begin
            S = 8'b00010000;
        end
    end
    if(A == 8'b00001001) begin
        if(B == 4'b1000) begin
            S = 8'b000010001;
        end
    end
    if(A == 8'b00001010) begin
        if(B == 4'b1000) begin
            S = 8'b000010010;
        end
    end
    if(A == 8'b00001011) begin
        if(B == 4'b1000) begin
            S = 8'b000010011;
        end
    end
    if(A == 8'b00001100) begin
        if(B == 4'b1000) begin
            S = 8'b000010100;
        end
    end
    if(A == 8'b00001101) begin
        if(B == 4'b1000) begin
            S = 8'b000010101;
        end
    end
    if(A == 8'b00001110) begin
        if(B == 4'b1000) begin
            S = 8'b000010110;
        end
    end
    if(A == 8'b00001111) begin
        if(B == 4'b1000) begin
            S = 8'b000010111;
        end
    end
    if(A == 8'b00010000) begin
        if(B == 4'b1000) begin
            S = 8'b00011000;
        end
    end
    if(A == 8'b000010001) begin
        if(B == 4'b1000) begin
            S = 8'b00011001;
        end
    end
    if(A == 8'b000010010) begin
        if(B == 4'b1000) begin
            S = 8'b00011010;
        end
    end
    if(A == 8'b000010011) begin
        if(B == 4'b1000) begin
            S = 8'b00011011;
        end
    end
    if(A == 8'b000010100) begin
        if(B == 4'b1000) begin
            S = 8'b00011100;
        end
    end
    if(A == 8'b000010101) begin
        if(B == 4'b1000) begin
            S = 8'b00011101;
        end
    end
    if(A == 8'b000010110) begin
        if(B == 4'b1000) begin
            S = 8'b00011110;
        end
    end
    if(A == 8'b000010111) begin
        if(B == 4'b1000) begin
            S = 8'b00011111;
        end
    end
    if(A == 8'b00011000) begin
        if(B == 4'b1000) begin
            S = 8'b00100000;
        end
    end
    if(A == 8'b00011001) begin
        if(B == 4'b1000) begin
            S = 8'b00100001;
        end
    end
    if(A == 8'b00011010) begin
        if(B == 4'b1000) begin
            S = 8'b00100010;
        end
    end
    if(A == 8'b00011011) begin
        if(B == 4'b1000) begin
            S = 8'b00100011;
        end
    end
    if(A == 8'b00011100) begin
        if(B == 4'b1000) begin
            S = 8'b00100100;
        end
    end
    if(A == 8'b00011101) begin
        if(B == 4'b1000) begin
            S = 8'b00100101;
        end
    end
    if(A == 8'b00011110) begin
        if(B == 4'b1000) begin
            S = 8'b00100110;
        end
    end
    if(A == 8'b00011111) begin
        if(B == 4'b1000) begin
            S = 8'b00100111;
        end
    end
    if(A == 8'b00100000) begin
        if(B == 4'b1000) begin
            S = 8'b00101000;
        end
    end
    if(A == 8'b00100001) begin
        if(B == 4'b1000) begin
            S = 8'b00101001;
        end
    end
    if(A == 8'b00100010) begin
        if(B == 4'b1000) begin
            S = 8'b00101010;
        end
    end
    if(A == 8'b00100011) begin
        if(B == 4'b1000) begin
            S = 8'b00101011;
        end
    end
    if(A == 8'b00100100) begin
        if(B == 4'b1000) begin
            S = 8'b00101100;
        end
    end
    if(A == 8'b00100101) begin
        if(B == 4'b1000) begin
            S = 8'b00101101;
        end
    end
    if(A == 8'b00100110) begin
        if(B == 4'b1000) begin
            S = 8'b00101110;
        end
    end
    if(A == 8'b00100111) begin
        if(B == 4'b1000) begin
            S = 8'b00101111;
        end
    end
    if(A == 8'b00101000) begin
        if(B == 4'b1000) begin
            S = 8'b00110000;
        end
    end
    if(A == 8'b00101001) begin
        if(B == 4'b1000) begin
            S = 8'b00110001;
        end
    end
    if(A == 8'b00101010) begin
        if(B == 4'b1000) begin
            S = 8'b00110010;
        end
    end
    if(A == 8'b00101011) begin
        if(B == 4'b1000) begin
            S = 8'b00110011;
        end
    end
    if(A == 8'b00101100) begin
        if(B == 4'b1000) begin
            S = 8'b00110100;
        end
    end
    if(A == 8'b00101101) begin
        if(B == 4'b1000) begin
            S = 8'b00110101;
        end
    end
    if(A == 8'b00101110) begin
        if(B == 4'b1000) begin
            S = 8'b00110110;
        end
    end
    if(A == 8'b00101111) begin
        if(B == 4'b1000) begin
            S = 8'b00110111;
        end
    end
    if(A == 8'b00110000) begin
        if(B == 4'b1000) begin
            S = 8'b00111000;
        end
    end
    if(A == 8'b00110001) begin
        if(B == 4'b1000) begin
            S = 8'b00111001;
        end
    end
    if(A == 8'b00110010) begin
        if(B == 4'b1000) begin
            S = 8'b00111010;
        end
    end
    if(A == 8'b00110011) begin
        if(B == 4'b1000) begin
            S = 8'b00111011;
        end
    end
    if(A == 8'b00110100) begin
        if(B == 4'b1000) begin
            S = 8'b00111100;
        end
    end
    if(A == 8'b00110101) begin
        if(B == 4'b1000) begin
            S = 8'b00111101;
        end
    end
    if(A == 8'b00110110) begin
        if(B == 4'b1000) begin
            S = 8'b00111110;
        end
    end
    if(A == 8'b00110111) begin
        if(B == 4'b1000) begin
            S = 8'b00111111;
        end
    end
    if(A == 8'b00111000) begin
        if(B == 4'b1000) begin
            S = 8'b01000000;
        end
    end
    if(A == 8'b00111001) begin
        if(B == 4'b1000) begin
            S = 8'b01000001;
        end
    end
    if(A == 8'b00111010) begin
        if(B == 4'b1000) begin
            S = 8'b01000010;
        end
    end
    if(A == 8'b00111011) begin
        if(B == 4'b1000) begin
            S = 8'b01000011;
        end
    end
    if(A == 8'b00111100) begin
        if(B == 4'b1000) begin
            S = 8'b01000100;
        end
    end
    if(A == 8'b00111101) begin
        if(B == 4'b1000) begin
            S = 8'b01000101;
        end
    end
    if(A == 8'b00111110) begin
        if(B == 4'b1000) begin
            S = 8'b01000110;
        end
    end
    if(A == 8'b00111111) begin
        if(B == 4'b1000) begin
            S = 8'b01000111;
        end
    end
    if(A == 8'b01000000) begin
        if(B == 4'b1000) begin
            S = 8'b01001000;
        end
    end
    if(A == 8'b01000001) begin
        if(B == 4'b1000) begin
            S = 8'b01001001;
        end
    end
    if(A == 8'b01000010) begin
        if(B == 4'b1000) begin
            S = 8'b01001010;
        end
    end
    if(A == 8'b01000011) begin
        if(B == 4'b1000) begin
            S = 8'b01001011;
        end
    end
    if(A == 8'b01000100) begin
        if(B == 4'b1000) begin
            S = 8'b01001100;
        end
    end
    if(A == 8'b01000101) begin
        if(B == 4'b1000) begin
            S = 8'b01001101;
        end
    end
    if(A == 8'b01000110) begin
        if(B == 4'b1000) begin
            S = 8'b01001110;
        end
    end
    if(A == 8'b01000111) begin
        if(B == 4'b1000) begin
            S = 8'b01001111;
        end
    end
    if(A == 8'b01001000) begin
        if(B == 4'b1000) begin
            S = 8'b01010000;
        end
    end
    if(A == 8'b01001001) begin
        if(B == 4'b1000) begin
            S = 8'b01010001;
        end
    end
    if(A == 8'b01001010) begin
        if(B == 4'b1000) begin
            S = 8'b01010010;
        end
    end
    if(A == 8'b01001011) begin
        if(B == 4'b1000) begin
            S = 8'b01010011;
        end
    end
    if(A == 8'b01001100) begin
        if(B == 4'b1000) begin
            S = 8'b01010100;
        end
    end
    if(A == 8'b01001101) begin
        if(B == 4'b1000) begin
            S = 8'b01010101;
        end
    end
    if(A == 8'b01001110) begin
        if(B == 4'b1000) begin
            S = 8'b01010110;
        end
    end
    if(A == 8'b01001111) begin
        if(B == 4'b1000) begin
            S = 8'b01010111;
        end
    end
    if(A == 8'b01010000) begin
        if(B == 4'b1000) begin
            S = 8'b01011000;
        end
    end
    if(A == 8'b01010001) begin
        if(B == 4'b1000) begin
            S = 8'b01011001;
        end
    end
    if(A == 8'b01010010) begin
        if(B == 4'b1000) begin
            S = 8'b01011010;
        end
    end
    if(A == 8'b01010011) begin
        if(B == 4'b1000) begin
            S = 8'b01011011;
        end
    end
    if(A == 8'b01010100) begin
        if(B == 4'b1000) begin
            S = 8'b01011100;
        end
    end
    if(A == 8'b01010101) begin
        if(B == 4'b1000) begin
            S = 8'b01011101;
        end
    end
    if(A == 8'b01010110) begin
        if(B == 4'b1000) begin
            S = 8'b01011110;
        end
    end
    if(A == 8'b01010111) begin
        if(B == 4'b1000) begin
            S = 8'b01011111;
        end
    end
    if(A == 8'b01011000) begin
        if(B == 4'b1000) begin
            S = 8'b01100000;
        end
    end
    if(A == 8'b01011001) begin
        if(B == 4'b1000) begin
            S = 8'b01100001;
        end
    end
    if(A == 8'b01011010) begin
        if(B == 4'b1000) begin
            S = 8'b01100010;
        end
    end
    if(A == 8'b01011011) begin
        if(B == 4'b1000) begin
            S = 8'b01100011;
        end
    end
    if(A == 8'b00000000) begin
        if(B == 4'b1001) begin
            S = 8'b00001001;
        end
    end
    if(A == 8'b00000001) begin
        if(B == 4'b1001) begin
            S = 8'b00001010;
        end
    end
    if(A == 8'b00000010) begin
        if(B == 4'b1001) begin
            S = 8'b00001011;
        end
    end
    if(A == 8'b00000011) begin
        if(B == 4'b1001) begin
            S = 8'b00001100;
        end
    end
    if(A == 8'b00000100) begin
        if(B == 4'b1001) begin
            S = 8'b00001101;
        end
    end
    if(A == 8'b00000101) begin
        if(B == 4'b1001) begin
            S = 8'b00001110;
        end
    end
    if(A == 8'b00000110) begin
        if(B == 4'b1001) begin
            S = 8'b00001111;
        end
    end
    if(A == 8'b00000111) begin
        if(B == 4'b1001) begin
            S = 8'b00010000;
        end
    end
    if(A == 8'b00001000) begin
        if(B == 4'b1001) begin
            S = 8'b000010001;
        end
    end
    if(A == 8'b00001001) begin
        if(B == 4'b1001) begin
            S = 8'b000010010;
        end
    end
    if(A == 8'b00001010) begin
        if(B == 4'b1001) begin
            S = 8'b000010011;
        end
    end
    if(A == 8'b00001011) begin
        if(B == 4'b1001) begin
            S = 8'b000010100;
        end
    end
    if(A == 8'b00001100) begin
        if(B == 4'b1001) begin
            S = 8'b000010101;
        end
    end
    if(A == 8'b00001101) begin
        if(B == 4'b1001) begin
            S = 8'b000010110;
        end
    end
    if(A == 8'b00001110) begin
        if(B == 4'b1001) begin
            S = 8'b000010111;
        end
    end
    if(A == 8'b00001111) begin
        if(B == 4'b1001) begin
            S = 8'b00011000;
        end
    end
    if(A == 8'b00010000) begin
        if(B == 4'b1001) begin
            S = 8'b00011001;
        end
    end
    if(A == 8'b000010001) begin
        if(B == 4'b1001) begin
            S = 8'b00011010;
        end
    end
    if(A == 8'b000010010) begin
        if(B == 4'b1001) begin
            S = 8'b00011011;
        end
    end
    if(A == 8'b000010011) begin
        if(B == 4'b1001) begin
            S = 8'b00011100;
        end
    end
    if(A == 8'b000010100) begin
        if(B == 4'b1001) begin
            S = 8'b00011101;
        end
    end
    if(A == 8'b000010101) begin
        if(B == 4'b1001) begin
            S = 8'b00011110;
        end
    end
    if(A == 8'b000010110) begin
        if(B == 4'b1001) begin
            S = 8'b00011111;
        end
    end
    if(A == 8'b000010111) begin
        if(B == 4'b1001) begin
            S = 8'b00100000;
        end
    end
    if(A == 8'b00011000) begin
        if(B == 4'b1001) begin
            S = 8'b00100001;
        end
    end
    if(A == 8'b00011001) begin
        if(B == 4'b1001) begin
            S = 8'b00100010;
        end
    end
    if(A == 8'b00011010) begin
        if(B == 4'b1001) begin
            S = 8'b00100011;
        end
    end
    if(A == 8'b00011011) begin
        if(B == 4'b1001) begin
            S = 8'b00100100;
        end
    end
    if(A == 8'b00011100) begin
        if(B == 4'b1001) begin
            S = 8'b00100101;
        end
    end
    if(A == 8'b00011101) begin
        if(B == 4'b1001) begin
            S = 8'b00100110;
        end
    end
    if(A == 8'b00011110) begin
        if(B == 4'b1001) begin
            S = 8'b00100111;
        end
    end
    if(A == 8'b00011111) begin
        if(B == 4'b1001) begin
            S = 8'b00101000;
        end
    end
    if(A == 8'b00100000) begin
        if(B == 4'b1001) begin
            S = 8'b00101001;
        end
    end
    if(A == 8'b00100001) begin
        if(B == 4'b1001) begin
            S = 8'b00101010;
        end
    end
    if(A == 8'b00100010) begin
        if(B == 4'b1001) begin
            S = 8'b00101011;
        end
    end
    if(A == 8'b00100011) begin
        if(B == 4'b1001) begin
            S = 8'b00101100;
        end
    end
    if(A == 8'b00100100) begin
        if(B == 4'b1001) begin
            S = 8'b00101101;
        end
    end
    if(A == 8'b00100101) begin
        if(B == 4'b1001) begin
            S = 8'b00101110;
        end
    end
    if(A == 8'b00100110) begin
        if(B == 4'b1001) begin
            S = 8'b00101111;
        end
    end
    if(A == 8'b00100111) begin
        if(B == 4'b1001) begin
            S = 8'b00110000;
        end
    end
    if(A == 8'b00101000) begin
        if(B == 4'b1001) begin
            S = 8'b00110001;
        end
    end
    if(A == 8'b00101001) begin
        if(B == 4'b1001) begin
            S = 8'b00110010;
        end
    end
    if(A == 8'b00101010) begin
        if(B == 4'b1001) begin
            S = 8'b00110011;
        end
    end
    if(A == 8'b00101011) begin
        if(B == 4'b1001) begin
            S = 8'b00110100;
        end
    end
    if(A == 8'b00101100) begin
        if(B == 4'b1001) begin
            S = 8'b00110101;
        end
    end
    if(A == 8'b00101101) begin
        if(B == 4'b1001) begin
            S = 8'b00110110;
        end
    end
    if(A == 8'b00101110) begin
        if(B == 4'b1001) begin
            S = 8'b00110111;
        end
    end
    if(A == 8'b00101111) begin
        if(B == 4'b1001) begin
            S = 8'b00111000;
        end
    end
    if(A == 8'b00110000) begin
        if(B == 4'b1001) begin
            S = 8'b00111001;
        end
    end
    if(A == 8'b00110001) begin
        if(B == 4'b1001) begin
            S = 8'b00111010;
        end
    end
    if(A == 8'b00110010) begin
        if(B == 4'b1001) begin
            S = 8'b00111011;
        end
    end
    if(A == 8'b00110011) begin
        if(B == 4'b1001) begin
            S = 8'b00111100;
        end
    end
    if(A == 8'b00110100) begin
        if(B == 4'b1001) begin
            S = 8'b00111101;
        end
    end
    if(A == 8'b00110101) begin
        if(B == 4'b1001) begin
            S = 8'b00111110;
        end
    end
    if(A == 8'b00110110) begin
        if(B == 4'b1001) begin
            S = 8'b00111111;
        end
    end
    if(A == 8'b00110111) begin
        if(B == 4'b1001) begin
            S = 8'b01000000;
        end
    end
    if(A == 8'b00111000) begin
        if(B == 4'b1001) begin
            S = 8'b01000001;
        end
    end
    if(A == 8'b00111001) begin
        if(B == 4'b1001) begin
            S = 8'b01000010;
        end
    end
    if(A == 8'b00111010) begin
        if(B == 4'b1001) begin
            S = 8'b01000011;
        end
    end
    if(A == 8'b00111011) begin
        if(B == 4'b1001) begin
            S = 8'b01000100;
        end
    end
    if(A == 8'b00111100) begin
        if(B == 4'b1001) begin
            S = 8'b01000101;
        end
    end
    if(A == 8'b00111101) begin
        if(B == 4'b1001) begin
            S = 8'b01000110;
        end
    end
    if(A == 8'b00111110) begin
        if(B == 4'b1001) begin
            S = 8'b01000111;
        end
    end
    if(A == 8'b00111111) begin
        if(B == 4'b1001) begin
            S = 8'b01001000;
        end
    end
    if(A == 8'b01000000) begin
        if(B == 4'b1001) begin
            S = 8'b01001001;
        end
    end
    if(A == 8'b01000001) begin
        if(B == 4'b1001) begin
            S = 8'b01001010;
        end
    end
    if(A == 8'b01000010) begin
        if(B == 4'b1001) begin
            S = 8'b01001011;
        end
    end
    if(A == 8'b01000011) begin
        if(B == 4'b1001) begin
            S = 8'b01001100;
        end
    end
    if(A == 8'b01000100) begin
        if(B == 4'b1001) begin
            S = 8'b01001101;
        end
    end
    if(A == 8'b01000101) begin
        if(B == 4'b1001) begin
            S = 8'b01001110;
        end
    end
    if(A == 8'b01000110) begin
        if(B == 4'b1001) begin
            S = 8'b01001111;
        end
    end
    if(A == 8'b01000111) begin
        if(B == 4'b1001) begin
            S = 8'b01010000;
        end
    end
    if(A == 8'b01001000) begin
        if(B == 4'b1001) begin
            S = 8'b01010001;
        end
    end
    if(A == 8'b01001001) begin
        if(B == 4'b1001) begin
            S = 8'b01010010;
        end
    end
    if(A == 8'b01001010) begin
        if(B == 4'b1001) begin
            S = 8'b01010011;
        end
    end
    if(A == 8'b01001011) begin
        if(B == 4'b1001) begin
            S = 8'b01010100;
        end
    end
    if(A == 8'b01001100) begin
        if(B == 4'b1001) begin
            S = 8'b01010101;
        end
    end
    if(A == 8'b01001101) begin
        if(B == 4'b1001) begin
            S = 8'b01010110;
        end
    end
    if(A == 8'b01001110) begin
        if(B == 4'b1001) begin
            S = 8'b01010111;
        end
    end
    if(A == 8'b01001111) begin
        if(B == 4'b1001) begin
            S = 8'b01011000;
        end
    end
    if(A == 8'b01010000) begin
        if(B == 4'b1001) begin
            S = 8'b01011001;
        end
    end
    if(A == 8'b01010001) begin
        if(B == 4'b1001) begin
            S = 8'b01011010;
        end
    end
    if(A == 8'b01010010) begin
        if(B == 4'b1001) begin
            S = 8'b01011011;
        end
    end
    if(A == 8'b01010011) begin
        if(B == 4'b1001) begin
            S = 8'b01011100;
        end
    end
    if(A == 8'b01010100) begin
        if(B == 4'b1001) begin
            S = 8'b01011101;
        end
    end
    if(A == 8'b01010101) begin
        if(B == 4'b1001) begin
            S = 8'b01011110;
        end
    end
    if(A == 8'b01010110) begin
        if(B == 4'b1001) begin
            S = 8'b01011111;
        end
    end
    if(A == 8'b01010111) begin
        if(B == 4'b1001) begin
            S = 8'b01100000;
        end
    end
    if(A == 8'b01011000) begin
        if(B == 4'b1001) begin
            S = 8'b01100001;
        end
    end
    if(A == 8'b01011001) begin
        if(B == 4'b1001) begin
            S = 8'b01100010;
        end
    end
    if(A == 8'b01011010) begin
        if(B == 4'b1001) begin
            S = 8'b01100011;
        end
    end
end
endmodule